`timescale 1 ps/ 1 ps

module ccgg(
	CI_CK,
	CI_CS,
	CI_DAT,
	CO_CK,
	CO_CS,
	CO_DAT,
	D0,
	D1,
	D10,
	D11,
	D12,
	D13,
	D14,
	D15,
	D16,
	D17,
	D18,
	D19,
	D2,
	D20,
	D21,
	D22,
	D23,
	D3,
	D4,
	D5,
	D6,
	D7,
	D8,
	D9,
	LM_CK,
	LM_D0,
	LM_D1,
	LM_D2,
	LM_D3,
	LM_D4,
	LM_D5,
	LM_LD,
	PIN_HSE,
	PIN_HSI,
	PIN_OSC,
	SH1,
	SH2,
	SH3,
	SH4,
	SH5,
	SH6,
	ST1,
	ST2);
input	CI_CK;
input	CI_CS;
input	CI_DAT;
output	CO_CK;
output	CO_CS;
output	CO_DAT;
output	D0;
output	D1;
output	D10;
output	D11;
output	D12;
output	D13;
output	D14;
output	D15;
output	D16;
output	D17;
output	D18;
output	D19;
output	D2;
output	D20;
output	D21;
output	D22;
output	D23;
output	D3;
output	D4;
output	D5;
output	D6;
output	D7;
output	D8;
output	D9;
output	LM_CK;
input	LM_D0;
input	LM_D1;
input	LM_D2;
input	LM_D3;
input	LM_D4;
input	LM_D5;
output	LM_LD;
input	PIN_HSE;
input	PIN_HSI;
input	PIN_OSC;
output	SH1;
output	SH2;
output	SH3;
output	SH4;
output	SH5;
output	SH6;
output	ST1;
output	ST2;

//wire	gnd;
//wire	vcc;
//wire	unknown;
wire	AsyncReset_X49_Y2_GND;
wire	AsyncReset_X49_Y3_GND;
wire	AsyncReset_X50_Y3_GND;
wire	AsyncReset_X51_Y3_GND;
wire	AsyncReset_X52_Y3_GND;
wire	\CI_CK~input_o ;
wire	\CI_CS~input_o ;
wire	\CI_DAT~input_o ;
wire	\LM_D0~input_o ;
wire	\LM_D1~input_o ;
wire	\LM_D2~input_o ;
wire	\LM_D3~input_o ;
wire	\LM_D4~input_o ;
wire	\LM_D5~input_o ;
wire	\PIN_HSE~input_o ;
wire	\PIN_HSI~input_o ;
wire	\PIN_OSC~input_o ;
wire	\PLL_ENABLE~clkctrl_outclk ;
wire	\PLL_ENABLE~clkctrl_outclk__AsyncReset_X48_Y1_SIG ;
wire	\PLL_ENABLE~combout ;
wire	\PLL_LOCK~combout ;
wire	SyncLoad_X43_Y2_GND;
wire	SyncLoad_X46_Y3_VCC;
wire	SyncLoad_X47_Y3_VCC;
wire	SyncLoad_X49_Y2_VCC;
wire	SyncLoad_X49_Y3_VCC;
wire	SyncLoad_X50_Y2_GND;
wire	SyncLoad_X50_Y3_VCC;
wire	SyncLoad_X51_Y2_GND;
wire	SyncLoad_X51_Y3_VCC;
wire	SyncLoad_X51_Y4_VCC;
wire	SyncLoad_X52_Y2_VCC;
wire	SyncLoad_X52_Y3_VCC;
wire	SyncLoad_X52_Y4_VCC;
wire	SyncLoad_X53_Y4_VCC;
wire	SyncLoad_X54_Y1_VCC;
wire	SyncLoad_X54_Y2_VCC;
wire	SyncLoad_X54_Y3_VCC;
wire	SyncLoad_X54_Y4_VCC;
wire	SyncLoad_X56_Y10_VCC;
wire	SyncLoad_X56_Y1_VCC;
wire	SyncLoad_X56_Y2_VCC;
wire	SyncLoad_X56_Y3_GND;
wire	SyncLoad_X56_Y4_VCC;
wire	SyncLoad_X56_Y5_GND;
wire	SyncLoad_X56_Y6_VCC;
wire	SyncLoad_X56_Y7_VCC;
wire	SyncLoad_X56_Y8_VCC;
wire	SyncLoad_X56_Y9_VCC;
wire	SyncLoad_X57_Y10_VCC;
wire	SyncLoad_X57_Y11_VCC;
wire	SyncLoad_X57_Y12_VCC;
wire	SyncLoad_X57_Y1_VCC;
wire	SyncLoad_X57_Y2_VCC;
wire	SyncLoad_X57_Y3_VCC;
wire	SyncLoad_X57_Y4_VCC;
wire	SyncLoad_X57_Y5_GND;
wire	SyncLoad_X57_Y6_VCC;
wire	SyncLoad_X57_Y8_VCC;
wire	SyncLoad_X57_Y9_VCC;
wire	SyncLoad_X58_Y10_VCC;
wire	SyncLoad_X58_Y11_VCC;
wire	SyncLoad_X58_Y12_VCC;
wire	SyncLoad_X58_Y1_VCC;
wire	SyncLoad_X58_Y2_VCC;
wire	SyncLoad_X58_Y3_VCC;
wire	SyncLoad_X58_Y4_VCC;
wire	SyncLoad_X58_Y5_VCC;
wire	SyncLoad_X58_Y6_VCC;
wire	SyncLoad_X58_Y7_VCC;
wire	SyncLoad_X58_Y8_VCC;
wire	SyncLoad_X58_Y9_VCC;
wire	SyncLoad_X59_Y10_VCC;
wire	SyncLoad_X59_Y11_VCC;
wire	SyncLoad_X59_Y12_VCC;
wire	SyncLoad_X59_Y1_VCC;
wire	SyncLoad_X59_Y2_VCC;
wire	SyncLoad_X59_Y3_VCC;
wire	SyncLoad_X59_Y4_VCC;
wire	SyncLoad_X59_Y5_VCC;
wire	SyncLoad_X59_Y7_VCC;
wire	SyncLoad_X59_Y8_VCC;
wire	SyncLoad_X59_Y9_VCC;
wire	SyncLoad_X60_Y10_VCC;
wire	SyncLoad_X60_Y11_VCC;
wire	SyncLoad_X60_Y12_VCC;
wire	SyncLoad_X60_Y1_VCC;
wire	SyncLoad_X60_Y2_VCC;
wire	SyncLoad_X60_Y3_VCC;
wire	SyncLoad_X60_Y4_VCC;
wire	SyncLoad_X60_Y5_VCC;
wire	SyncLoad_X60_Y6_VCC;
wire	SyncLoad_X60_Y7_VCC;
wire	SyncLoad_X60_Y8_VCC;
wire	SyncLoad_X60_Y9_VCC;
wire	SyncLoad_X61_Y10_VCC;
wire	SyncLoad_X61_Y11_VCC;
wire	SyncLoad_X61_Y1_VCC;
wire	SyncLoad_X61_Y2_VCC;
wire	SyncLoad_X61_Y3_VCC;
wire	SyncLoad_X61_Y4_VCC;
wire	SyncLoad_X61_Y5_VCC;
wire	SyncLoad_X61_Y6_VCC;
wire	SyncLoad_X61_Y7_VCC;
wire	SyncLoad_X61_Y8_VCC;
wire	SyncLoad_X61_Y9_VCC;
wire	SyncLoad_X62_Y10_VCC;
wire	SyncLoad_X62_Y11_VCC;
wire	SyncLoad_X62_Y1_VCC;
wire	SyncLoad_X62_Y2_VCC;
wire	SyncLoad_X62_Y3_VCC;
wire	SyncLoad_X62_Y4_VCC;
wire	SyncLoad_X62_Y5_VCC;
wire	SyncLoad_X62_Y6_VCC;
wire	SyncLoad_X62_Y7_VCC;
wire	SyncLoad_X62_Y8_VCC;
wire	SyncLoad_X62_Y9_VCC;
wire	SyncReset_X46_Y2_GND;
wire	SyncReset_X46_Y3_GND;
wire	SyncReset_X47_Y3_GND;
wire	SyncReset_X49_Y2_GND;
wire	SyncReset_X49_Y3_GND;
wire	SyncReset_X50_Y1_GND;
wire	SyncReset_X50_Y3_GND;
wire	SyncReset_X51_Y3_GND;
wire	SyncReset_X51_Y4_GND;
wire	SyncReset_X52_Y2_GND;
wire	SyncReset_X52_Y3_GND;
wire	SyncReset_X52_Y4_GND;
wire	SyncReset_X53_Y4_GND;
wire	SyncReset_X54_Y1_GND;
wire	SyncReset_X54_Y2_GND;
wire	SyncReset_X54_Y3_GND;
wire	SyncReset_X54_Y4_GND;
wire	SyncReset_X56_Y10_GND;
wire	SyncReset_X56_Y1_GND;
wire	SyncReset_X56_Y2_GND;
wire	SyncReset_X56_Y4_GND;
wire	SyncReset_X56_Y6_GND;
wire	SyncReset_X56_Y7_GND;
wire	SyncReset_X56_Y8_GND;
wire	SyncReset_X56_Y9_GND;
wire	SyncReset_X57_Y10_GND;
wire	SyncReset_X57_Y11_GND;
wire	SyncReset_X57_Y12_GND;
wire	SyncReset_X57_Y1_GND;
wire	SyncReset_X57_Y2_GND;
wire	SyncReset_X57_Y3_GND;
wire	SyncReset_X57_Y4_GND;
wire	SyncReset_X57_Y6_GND;
wire	SyncReset_X57_Y8_GND;
wire	SyncReset_X57_Y9_GND;
wire	SyncReset_X58_Y10_GND;
wire	SyncReset_X58_Y11_GND;
wire	SyncReset_X58_Y12_GND;
wire	SyncReset_X58_Y1_GND;
wire	SyncReset_X58_Y2_GND;
wire	SyncReset_X58_Y3_GND;
wire	SyncReset_X58_Y4_GND;
wire	SyncReset_X58_Y5_GND;
wire	SyncReset_X58_Y6_GND;
wire	SyncReset_X58_Y7_GND;
wire	SyncReset_X58_Y8_GND;
wire	SyncReset_X58_Y9_GND;
wire	SyncReset_X59_Y10_GND;
wire	SyncReset_X59_Y11_GND;
wire	SyncReset_X59_Y12_GND;
wire	SyncReset_X59_Y1_GND;
wire	SyncReset_X59_Y2_GND;
wire	SyncReset_X59_Y3_GND;
wire	SyncReset_X59_Y4_GND;
wire	SyncReset_X59_Y5_GND;
wire	SyncReset_X59_Y7_GND;
wire	SyncReset_X59_Y8_GND;
wire	SyncReset_X59_Y9_GND;
wire	SyncReset_X60_Y10_GND;
wire	SyncReset_X60_Y11_GND;
wire	SyncReset_X60_Y12_GND;
wire	SyncReset_X60_Y1_GND;
wire	SyncReset_X60_Y2_GND;
wire	SyncReset_X60_Y3_GND;
wire	SyncReset_X60_Y4_GND;
wire	SyncReset_X60_Y5_GND;
wire	SyncReset_X60_Y6_GND;
wire	SyncReset_X60_Y7_GND;
wire	SyncReset_X60_Y8_GND;
wire	SyncReset_X60_Y9_GND;
wire	SyncReset_X61_Y10_GND;
wire	SyncReset_X61_Y11_GND;
wire	SyncReset_X61_Y1_GND;
wire	SyncReset_X61_Y2_GND;
wire	SyncReset_X61_Y3_GND;
wire	SyncReset_X61_Y4_GND;
wire	SyncReset_X61_Y5_GND;
wire	SyncReset_X61_Y6_GND;
wire	SyncReset_X61_Y7_GND;
wire	SyncReset_X61_Y8_GND;
wire	SyncReset_X61_Y9_GND;
wire	SyncReset_X62_Y10_GND;
wire	SyncReset_X62_Y11_GND;
wire	SyncReset_X62_Y1_GND;
wire	SyncReset_X62_Y2_GND;
wire	SyncReset_X62_Y3_GND;
wire	SyncReset_X62_Y4_GND;
wire	SyncReset_X62_Y5_GND;
wire	SyncReset_X62_Y6_GND;
wire	SyncReset_X62_Y7_GND;
wire	SyncReset_X62_Y8_GND;
wire	SyncReset_X62_Y9_GND;
wire	\auto_generated_inst.hbo_13_1bc039b416d3bc4a_bp ;
wire	\auto_generated_inst.hbo_13_1bc039b416d3bc4a_bp_X48_Y1_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X46_Y3_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X47_Y2_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X47_Y3_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y2_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y3_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X49_Y1_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X49_Y4_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X50_Y1_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X51_Y1_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X54_Y2_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X54_Y4_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y10_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y11_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y1_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y4_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y6_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y7_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y9_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y12_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y1_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y2_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y3_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y4_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y7_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y9_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y11_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y12_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y4_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y7_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y10_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y12_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y1_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y2_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y3_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y5_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X60_Y1_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X60_Y6_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y11_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y12_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y2_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y5_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y8_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y9_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y10_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y12_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y1_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y3_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y4_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y5_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y7_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y8_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y9_SIG_VCC ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X54_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X57_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X58_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X59_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X60_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|pwmUpdateTrigger~q_X59_Y6_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|Equal0~0_combout_X50_Y1_SIG_INV ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|bit_counter[7]~8_combout_X50_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|byte_counter[4]~10_combout_X51_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|scaler_counter[0]~0_combout_X51_Y1_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X51_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X52_Y1_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X52_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X53_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X50_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y11_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X59_Y8_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y1_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y11_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X59_Y7_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X60_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X57_Y6_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X58_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X58_Y5_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X59_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X56_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X57_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X61_Y6_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X62_Y6_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X57_Y8_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y8_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y9_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X58_Y5_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X60_Y5_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X57_Y11_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X59_Y9_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X59_Y12_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X60_Y12_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X57_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X58_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X60_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X61_Y5_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X56_Y8_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X62_Y8_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X59_Y11_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X60_Y11_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X60_Y6_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X61_Y10_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X59_Y10_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X60_Y12_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X57_Y6_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X57_Y7_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X58_Y10_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X60_Y1_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X61_Y1_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X58_Y10_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X60_Y8_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X62_Y6_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X58_Y12_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X59_Y11_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X60_Y9_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X58_Y6_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X61_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X62_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X58_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y8_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X60_Y7_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X61_Y7_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X60_Y8_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X62_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X59_Y6_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X59_Y9_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X60_Y7_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X61_Y11_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X56_Y10_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X57_Y10_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X54_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X60_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X56_Y1_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X58_Y1_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X56_Y9_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X58_Y9_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X56_Y6_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X60_Y10_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y7_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y8_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X57_Y9_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X60_Y5_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X60_Y9_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X61_Y9_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X56_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X59_Y7_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X57_Y8_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X58_Y7_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X61_Y6_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X62_Y5_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y10_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y12_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X58_Y8_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X60_Y10_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X62_Y9_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y11_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y7_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X59_Y5_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X60_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X57_Y1_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X58_Y1_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X58_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X59_Y1_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X60_Y11_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X61_Y8_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X61_Y10_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X62_Y10_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X57_Y11_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X58_Y11_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X61_Y7_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X62_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X56_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X59_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X54_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X58_Y6_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X60_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X61_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X62_Y1_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~1_combout_X50_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~2_combout_X51_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~3_combout_X52_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~4_combout_X49_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~5_combout_X49_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~6_combout_X52_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~7_combout_X49_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~8_combout_X50_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X54_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y5_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X57_Y5_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X49_Y2_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X49_Y4_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X51_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y3_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y5_SIG_SIG ;
wire	\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ;
tri1	devclrn;
tri1	devoe;
tri1	devpor;
wire	\gclksw_inst|gclk_switch__alta_gclksw__clkout ;
wire	hbi_272_0_9cb2c0024f9919c5_bp;
wire	hbi_272_1_9cb2c0024f9919c5_bp;
wire	\macro_inst|Add0~0_combout ;
wire	\macro_inst|Add0~1 ;
wire	\macro_inst|Add0~10_combout ;
wire	\macro_inst|Add0~11 ;
wire	\macro_inst|Add0~12_combout ;
wire	\macro_inst|Add0~13 ;
wire	\macro_inst|Add0~14_combout ;
wire	\macro_inst|Add0~15 ;
wire	\macro_inst|Add0~16_combout ;
wire	\macro_inst|Add0~17 ;
wire	\macro_inst|Add0~18_combout ;
wire	\macro_inst|Add0~19 ;
wire	\macro_inst|Add0~20_combout ;
wire	\macro_inst|Add0~21 ;
wire	\macro_inst|Add0~22_combout ;
wire	\macro_inst|Add0~23 ;
wire	\macro_inst|Add0~24_combout ;
wire	\macro_inst|Add0~25 ;
wire	\macro_inst|Add0~26_combout ;
wire	\macro_inst|Add0~27 ;
wire	\macro_inst|Add0~28_combout ;
wire	\macro_inst|Add0~29 ;
wire	\macro_inst|Add0~2_combout ;
wire	\macro_inst|Add0~3 ;
wire	\macro_inst|Add0~30_combout ;
wire	\macro_inst|Add0~31 ;
wire	\macro_inst|Add0~32_combout ;
wire	\macro_inst|Add0~33 ;
wire	\macro_inst|Add0~34_combout ;
wire	\macro_inst|Add0~35 ;
wire	\macro_inst|Add0~36_combout ;
wire	\macro_inst|Add0~37 ;
wire	\macro_inst|Add0~38_combout ;
wire	\macro_inst|Add0~39 ;
wire	\macro_inst|Add0~40_combout ;
wire	\macro_inst|Add0~41 ;
wire	\macro_inst|Add0~42_combout ;
wire	\macro_inst|Add0~43 ;
wire	\macro_inst|Add0~44_combout ;
wire	\macro_inst|Add0~4_combout ;
wire	\macro_inst|Add0~5 ;
wire	\macro_inst|Add0~6_combout ;
wire	\macro_inst|Add0~7 ;
wire	\macro_inst|Add0~8_combout ;
wire	\macro_inst|Add0~9 ;
wire	\macro_inst|Equal1~0_combout ;
wire	\macro_inst|Equal1~1_combout ;
wire	\macro_inst|Equal1~2_combout ;
wire	\macro_inst|Equal1~3_combout ;
wire	\macro_inst|Equal1~4_combout ;
wire	\macro_inst|Equal1~5_combout ;
wire	\macro_inst|Equal1~6_combout ;
wire	\macro_inst|Equal1~7_combout ;
wire	\macro_inst|Equal1~8_combout ;
wire	\macro_inst|Equal2~0_combout ;
wire	\macro_inst|Equal3~0_combout ;
wire	\macro_inst|Equal3~1_combout ;
wire	\macro_inst|Equal3~2_combout ;
wire	\macro_inst|Equal3~3_combout ;
wire	\macro_inst|Equal3~4_combout ;
wire	\macro_inst|Equal3~5_combout ;
wire	\macro_inst|Equal3~6_combout ;
wire	[31:0] \macro_inst|ahb_add_reg ;
//wire	\macro_inst|ahb_add_reg [0];
//wire	\macro_inst|ahb_add_reg [10];
//wire	\macro_inst|ahb_add_reg [11];
//wire	\macro_inst|ahb_add_reg [12];
//wire	\macro_inst|ahb_add_reg [13];
//wire	\macro_inst|ahb_add_reg [14];
//wire	\macro_inst|ahb_add_reg [15];
//wire	\macro_inst|ahb_add_reg [16];
//wire	\macro_inst|ahb_add_reg [17];
//wire	\macro_inst|ahb_add_reg [18];
//wire	\macro_inst|ahb_add_reg [19];
//wire	\macro_inst|ahb_add_reg [1];
//wire	\macro_inst|ahb_add_reg [20];
//wire	\macro_inst|ahb_add_reg [21];
//wire	\macro_inst|ahb_add_reg [22];
//wire	\macro_inst|ahb_add_reg [23];
//wire	\macro_inst|ahb_add_reg [24];
//wire	\macro_inst|ahb_add_reg [25];
//wire	\macro_inst|ahb_add_reg [26];
//wire	\macro_inst|ahb_add_reg [27];
//wire	\macro_inst|ahb_add_reg [28];
//wire	\macro_inst|ahb_add_reg [29];
//wire	\macro_inst|ahb_add_reg [2];
//wire	\macro_inst|ahb_add_reg [30];
//wire	\macro_inst|ahb_add_reg [31];
//wire	\macro_inst|ahb_add_reg [3];
//wire	\macro_inst|ahb_add_reg [4];
//wire	\macro_inst|ahb_add_reg [5];
//wire	\macro_inst|ahb_add_reg [6];
//wire	\macro_inst|ahb_add_reg [7];
//wire	\macro_inst|ahb_add_reg [8];
//wire	\macro_inst|ahb_add_reg [9];
wire	\macro_inst|ahb_ready_reg~q ;
wire	\macro_inst|ahb_wr_reg~q ;
wire	[22:0] \macro_inst|clk10hz_cnt ;
//wire	\macro_inst|clk10hz_cnt [0];
//wire	\macro_inst|clk10hz_cnt [10];
//wire	\macro_inst|clk10hz_cnt [11];
//wire	\macro_inst|clk10hz_cnt [12];
//wire	\macro_inst|clk10hz_cnt [13];
//wire	\macro_inst|clk10hz_cnt [14];
//wire	\macro_inst|clk10hz_cnt [15];
//wire	\macro_inst|clk10hz_cnt [16];
//wire	\macro_inst|clk10hz_cnt [17];
//wire	\macro_inst|clk10hz_cnt [18];
//wire	\macro_inst|clk10hz_cnt [19];
//wire	\macro_inst|clk10hz_cnt [1];
//wire	\macro_inst|clk10hz_cnt [20];
//wire	\macro_inst|clk10hz_cnt [21];
//wire	\macro_inst|clk10hz_cnt [22];
//wire	\macro_inst|clk10hz_cnt [2];
//wire	\macro_inst|clk10hz_cnt [3];
//wire	\macro_inst|clk10hz_cnt [4];
//wire	\macro_inst|clk10hz_cnt [5];
//wire	\macro_inst|clk10hz_cnt [6];
//wire	\macro_inst|clk10hz_cnt [7];
//wire	\macro_inst|clk10hz_cnt [8];
//wire	\macro_inst|clk10hz_cnt [9];
wire	\macro_inst|clk10hz_cnt~0_combout ;
wire	\macro_inst|clk10hz_cnt~1_combout ;
wire	\macro_inst|clk10hz_cnt~2_combout ;
wire	\macro_inst|clk10hz_cnt~3_combout ;
wire	\macro_inst|clk10hz_cnt~4_combout ;
wire	\macro_inst|clk10hz_cnt~5_combout ;
wire	\macro_inst|clock10Hz~0_combout ;
wire	\macro_inst|clock10Hz~q ;
wire	\macro_inst|controller|Add0~0_combout ;
wire	\macro_inst|controller|Add0~1 ;
wire	\macro_inst|controller|Add0~10_combout ;
wire	\macro_inst|controller|Add0~11 ;
wire	\macro_inst|controller|Add0~12_combout ;
wire	\macro_inst|controller|Add0~13 ;
wire	\macro_inst|controller|Add0~14_combout ;
wire	\macro_inst|controller|Add0~2_combout ;
wire	\macro_inst|controller|Add0~3 ;
wire	\macro_inst|controller|Add0~4_combout ;
wire	\macro_inst|controller|Add0~5 ;
wire	\macro_inst|controller|Add0~6_combout ;
wire	\macro_inst|controller|Add0~7 ;
wire	\macro_inst|controller|Add0~8_combout ;
wire	\macro_inst|controller|Add0~9 ;
wire	\macro_inst|controller|Equal1~0_combout ;
wire	\macro_inst|controller|Equal1~1_combout ;
wire	\macro_inst|controller|Equal1~2_combout ;
wire	\macro_inst|controller|pwmUpdateTrigger~feeder_combout ;
wire	\macro_inst|controller|pwmUpdateTrigger~q ;
wire	[1:0] \macro_inst|controller|serialOutputTrigger ;
//wire	\macro_inst|controller|serialOutputTrigger [0];
wire	\macro_inst|controller|serialOutputTrigger[0]~1_combout ;
//wire	\macro_inst|controller|serialOutputTrigger [1];
wire	\macro_inst|controller|serialOutputTrigger[1]~0_combout ;
wire	[7:0] \macro_inst|controller|serialTrigCounter ;
//wire	\macro_inst|controller|serialTrigCounter [0];
//wire	\macro_inst|controller|serialTrigCounter [1];
//wire	\macro_inst|controller|serialTrigCounter [2];
//wire	\macro_inst|controller|serialTrigCounter [3];
//wire	\macro_inst|controller|serialTrigCounter [4];
//wire	\macro_inst|controller|serialTrigCounter [5];
//wire	\macro_inst|controller|serialTrigCounter [6];
//wire	\macro_inst|controller|serialTrigCounter [7];
wire	\macro_inst|controller|serialTrigCounter~0_combout ;
wire	\macro_inst|controller|serialTrigCounter~1_combout ;
wire	\macro_inst|controller|serialTrigCounter~2_combout ;
wire	\macro_inst|controller|serial|Add2~0_combout ;
wire	\macro_inst|controller|serial|Add2~1_combout ;
wire	\macro_inst|controller|serial|Equal0~0_combout ;
wire	\macro_inst|controller|serial|Equal1~0_combout ;
wire	\macro_inst|controller|serial|Equal1~1_combout ;
wire	\macro_inst|controller|serial|Selector2~0_combout ;
wire	\macro_inst|controller|serial|Selector4~0_combout ;
wire	\macro_inst|controller|serial|Selector4~1_combout ;
wire	\macro_inst|controller|serial|Selector4~2_combout ;
wire	\macro_inst|controller|serial|Selector4~3_combout ;
wire	[7:0] \macro_inst|controller|serial|bit_counter ;
//wire	\macro_inst|controller|serial|bit_counter [0];
wire	\macro_inst|controller|serial|bit_counter[0]~10 ;
wire	\macro_inst|controller|serial|bit_counter[0]~9_combout ;
//wire	\macro_inst|controller|serial|bit_counter [1];
wire	\macro_inst|controller|serial|bit_counter[1]~11_combout ;
wire	\macro_inst|controller|serial|bit_counter[1]~12 ;
//wire	\macro_inst|controller|serial|bit_counter [2];
wire	\macro_inst|controller|serial|bit_counter[2]~13_combout ;
wire	\macro_inst|controller|serial|bit_counter[2]~14 ;
//wire	\macro_inst|controller|serial|bit_counter [3];
wire	\macro_inst|controller|serial|bit_counter[3]~15_combout ;
wire	\macro_inst|controller|serial|bit_counter[3]~16 ;
//wire	\macro_inst|controller|serial|bit_counter [4];
wire	\macro_inst|controller|serial|bit_counter[4]~18_combout ;
wire	\macro_inst|controller|serial|bit_counter[4]~19 ;
//wire	\macro_inst|controller|serial|bit_counter [5];
wire	\macro_inst|controller|serial|bit_counter[5]~20_combout ;
wire	\macro_inst|controller|serial|bit_counter[5]~21 ;
//wire	\macro_inst|controller|serial|bit_counter [6];
wire	\macro_inst|controller|serial|bit_counter[6]~22_combout ;
wire	\macro_inst|controller|serial|bit_counter[6]~23 ;
//wire	\macro_inst|controller|serial|bit_counter [7];
wire	\macro_inst|controller|serial|bit_counter[7]~17_combout ;
wire	\macro_inst|controller|serial|bit_counter[7]~17_combout__SyncReset_X50_Y2_SIG ;
wire	\macro_inst|controller|serial|bit_counter[7]~24_combout ;
wire	\macro_inst|controller|serial|bit_counter[7]~8_combout ;
wire	[7:0] \macro_inst|controller|serial|byte_counter ;
//wire	\macro_inst|controller|serial|byte_counter [0];
wire	\macro_inst|controller|serial|byte_counter[0]~8_combout ;
wire	\macro_inst|controller|serial|byte_counter[0]~9 ;
//wire	\macro_inst|controller|serial|byte_counter [1];
wire	\macro_inst|controller|serial|byte_counter[1]~11_combout ;
wire	\macro_inst|controller|serial|byte_counter[1]~12 ;
//wire	\macro_inst|controller|serial|byte_counter [2];
wire	\macro_inst|controller|serial|byte_counter[2]~13_combout ;
wire	\macro_inst|controller|serial|byte_counter[2]~14 ;
//wire	\macro_inst|controller|serial|byte_counter [3];
wire	\macro_inst|controller|serial|byte_counter[3]~15_combout ;
wire	\macro_inst|controller|serial|byte_counter[3]~16 ;
//wire	\macro_inst|controller|serial|byte_counter [4];
wire	\macro_inst|controller|serial|byte_counter[4]~10_combout ;
wire	\macro_inst|controller|serial|byte_counter[4]~17_combout ;
wire	\macro_inst|controller|serial|byte_counter[4]~18 ;
//wire	\macro_inst|controller|serial|byte_counter [5];
wire	\macro_inst|controller|serial|byte_counter[5]~19_combout ;
wire	\macro_inst|controller|serial|byte_counter[5]~20 ;
//wire	\macro_inst|controller|serial|byte_counter [6];
wire	\macro_inst|controller|serial|byte_counter[6]~21_combout ;
wire	\macro_inst|controller|serial|byte_counter[6]~22 ;
//wire	\macro_inst|controller|serial|byte_counter [7];
wire	\macro_inst|controller|serial|byte_counter[7]~23_combout ;
wire	[3:0] \macro_inst|controller|serial|scaler_counter ;
//wire	\macro_inst|controller|serial|scaler_counter [0];
wire	\macro_inst|controller|serial|scaler_counter[0]~0_combout ;
//wire	\macro_inst|controller|serial|scaler_counter [1];
//wire	\macro_inst|controller|serial|scaler_counter [2];
//wire	\macro_inst|controller|serial|scaler_counter [3];
wire	\macro_inst|controller|serial|scaler_counter~1_combout ;
wire	\macro_inst|controller|serial|scaler_counter~2_combout ;
wire	\macro_inst|controller|serial|scaler_counter~3_combout ;
wire	\macro_inst|controller|serial|scaler_counter~4_combout ;
wire	[23:0] \macro_inst|controller|serial|sdata_reg ;
//wire	\macro_inst|controller|serial|sdata_reg [0];
wire	\macro_inst|controller|serial|sdata_reg[0]~0_combout ;
wire	\macro_inst|controller|serial|sdata_reg[0]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [10];
wire	\macro_inst|controller|serial|sdata_reg[10]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [11];
wire	\macro_inst|controller|serial|sdata_reg[11]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [12];
//wire	\macro_inst|controller|serial|sdata_reg [13];
wire	\macro_inst|controller|serial|sdata_reg[13]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [14];
//wire	\macro_inst|controller|serial|sdata_reg [15];
wire	\macro_inst|controller|serial|sdata_reg[15]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [16];
wire	\macro_inst|controller|serial|sdata_reg[16]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [17];
wire	\macro_inst|controller|serial|sdata_reg[17]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [18];
wire	\macro_inst|controller|serial|sdata_reg[18]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [19];
wire	\macro_inst|controller|serial|sdata_reg[19]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [1];
wire	\macro_inst|controller|serial|sdata_reg[1]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [20];
//wire	\macro_inst|controller|serial|sdata_reg [21];
wire	\macro_inst|controller|serial|sdata_reg[21]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [22];
//wire	\macro_inst|controller|serial|sdata_reg [23];
//wire	\macro_inst|controller|serial|sdata_reg [2];
wire	\macro_inst|controller|serial|sdata_reg[2]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [3];
wire	\macro_inst|controller|serial|sdata_reg[3]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [4];
//wire	\macro_inst|controller|serial|sdata_reg [5];
wire	\macro_inst|controller|serial|sdata_reg[5]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [6];
wire	\macro_inst|controller|serial|sdata_reg[6]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [7];
wire	\macro_inst|controller|serial|sdata_reg[7]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [8];
wire	\macro_inst|controller|serial|sdata_reg[8]~feeder_combout ;
//wire	\macro_inst|controller|serial|sdata_reg [9];
wire	\macro_inst|controller|serial|sdata_reg[9]~feeder_combout ;
wire	[191:0] \macro_inst|controller|serial|shift_data ;
//wire	\macro_inst|controller|serial|shift_data [0];
//wire	\macro_inst|controller|serial|shift_data [100];
//wire	\macro_inst|controller|serial|shift_data [101];
//wire	\macro_inst|controller|serial|shift_data [102];
//wire	\macro_inst|controller|serial|shift_data [103];
//wire	\macro_inst|controller|serial|shift_data [104];
//wire	\macro_inst|controller|serial|shift_data [105];
//wire	\macro_inst|controller|serial|shift_data [106];
//wire	\macro_inst|controller|serial|shift_data [107];
//wire	\macro_inst|controller|serial|shift_data [108];
//wire	\macro_inst|controller|serial|shift_data [109];
//wire	\macro_inst|controller|serial|shift_data [10];
//wire	\macro_inst|controller|serial|shift_data [110];
//wire	\macro_inst|controller|serial|shift_data [111];
//wire	\macro_inst|controller|serial|shift_data [112];
//wire	\macro_inst|controller|serial|shift_data [113];
//wire	\macro_inst|controller|serial|shift_data [114];
//wire	\macro_inst|controller|serial|shift_data [115];
//wire	\macro_inst|controller|serial|shift_data [116];
//wire	\macro_inst|controller|serial|shift_data [117];
//wire	\macro_inst|controller|serial|shift_data [118];
//wire	\macro_inst|controller|serial|shift_data [119];
//wire	\macro_inst|controller|serial|shift_data [11];
//wire	\macro_inst|controller|serial|shift_data [120];
//wire	\macro_inst|controller|serial|shift_data [121];
//wire	\macro_inst|controller|serial|shift_data [122];
//wire	\macro_inst|controller|serial|shift_data [123];
//wire	\macro_inst|controller|serial|shift_data [124];
//wire	\macro_inst|controller|serial|shift_data [125];
//wire	\macro_inst|controller|serial|shift_data [126];
//wire	\macro_inst|controller|serial|shift_data [127];
//wire	\macro_inst|controller|serial|shift_data [128];
//wire	\macro_inst|controller|serial|shift_data [129];
//wire	\macro_inst|controller|serial|shift_data [12];
//wire	\macro_inst|controller|serial|shift_data [130];
//wire	\macro_inst|controller|serial|shift_data [131];
//wire	\macro_inst|controller|serial|shift_data [132];
//wire	\macro_inst|controller|serial|shift_data [133];
wire	\macro_inst|controller|serial|shift_data[133]~feeder_combout ;
//wire	\macro_inst|controller|serial|shift_data [134];
//wire	\macro_inst|controller|serial|shift_data [135];
//wire	\macro_inst|controller|serial|shift_data [136];
//wire	\macro_inst|controller|serial|shift_data [137];
//wire	\macro_inst|controller|serial|shift_data [138];
//wire	\macro_inst|controller|serial|shift_data [139];
//wire	\macro_inst|controller|serial|shift_data [13];
//wire	\macro_inst|controller|serial|shift_data [140];
//wire	\macro_inst|controller|serial|shift_data [141];
//wire	\macro_inst|controller|serial|shift_data [142];
//wire	\macro_inst|controller|serial|shift_data [143];
//wire	\macro_inst|controller|serial|shift_data [144];
//wire	\macro_inst|controller|serial|shift_data [145];
//wire	\macro_inst|controller|serial|shift_data [146];
//wire	\macro_inst|controller|serial|shift_data [147];
//wire	\macro_inst|controller|serial|shift_data [148];
//wire	\macro_inst|controller|serial|shift_data [149];
//wire	\macro_inst|controller|serial|shift_data [14];
//wire	\macro_inst|controller|serial|shift_data [150];
//wire	\macro_inst|controller|serial|shift_data [151];
//wire	\macro_inst|controller|serial|shift_data [152];
//wire	\macro_inst|controller|serial|shift_data [153];
//wire	\macro_inst|controller|serial|shift_data [154];
//wire	\macro_inst|controller|serial|shift_data [155];
//wire	\macro_inst|controller|serial|shift_data [156];
//wire	\macro_inst|controller|serial|shift_data [157];
//wire	\macro_inst|controller|serial|shift_data [158];
//wire	\macro_inst|controller|serial|shift_data [159];
//wire	\macro_inst|controller|serial|shift_data [15];
//wire	\macro_inst|controller|serial|shift_data [160];
//wire	\macro_inst|controller|serial|shift_data [161];
//wire	\macro_inst|controller|serial|shift_data [162];
//wire	\macro_inst|controller|serial|shift_data [163];
//wire	\macro_inst|controller|serial|shift_data [164];
//wire	\macro_inst|controller|serial|shift_data [165];
//wire	\macro_inst|controller|serial|shift_data [166];
//wire	\macro_inst|controller|serial|shift_data [167];
//wire	\macro_inst|controller|serial|shift_data [168];
//wire	\macro_inst|controller|serial|shift_data [169];
//wire	\macro_inst|controller|serial|shift_data [16];
//wire	\macro_inst|controller|serial|shift_data [170];
//wire	\macro_inst|controller|serial|shift_data [171];
//wire	\macro_inst|controller|serial|shift_data [172];
//wire	\macro_inst|controller|serial|shift_data [173];
//wire	\macro_inst|controller|serial|shift_data [174];
//wire	\macro_inst|controller|serial|shift_data [175];
//wire	\macro_inst|controller|serial|shift_data [176];
//wire	\macro_inst|controller|serial|shift_data [177];
//wire	\macro_inst|controller|serial|shift_data [178];
//wire	\macro_inst|controller|serial|shift_data [179];
//wire	\macro_inst|controller|serial|shift_data [17];
//wire	\macro_inst|controller|serial|shift_data [180];
//wire	\macro_inst|controller|serial|shift_data [181];
//wire	\macro_inst|controller|serial|shift_data [182];
//wire	\macro_inst|controller|serial|shift_data [183];
//wire	\macro_inst|controller|serial|shift_data [184];
//wire	\macro_inst|controller|serial|shift_data [185];
wire	\macro_inst|controller|serial|shift_data[185]~feeder_combout ;
//wire	\macro_inst|controller|serial|shift_data [186];
wire	\macro_inst|controller|serial|shift_data[186]~feeder_combout ;
//wire	\macro_inst|controller|serial|shift_data [187];
//wire	\macro_inst|controller|serial|shift_data [188];
//wire	\macro_inst|controller|serial|shift_data [189];
//wire	\macro_inst|controller|serial|shift_data [18];
//wire	\macro_inst|controller|serial|shift_data [190];
//wire	\macro_inst|controller|serial|shift_data [191];
//wire	\macro_inst|controller|serial|shift_data [19];
//wire	\macro_inst|controller|serial|shift_data [1];
//wire	\macro_inst|controller|serial|shift_data [20];
//wire	\macro_inst|controller|serial|shift_data [21];
//wire	\macro_inst|controller|serial|shift_data [22];
//wire	\macro_inst|controller|serial|shift_data [23];
//wire	\macro_inst|controller|serial|shift_data [24];
//wire	\macro_inst|controller|serial|shift_data [25];
//wire	\macro_inst|controller|serial|shift_data [26];
//wire	\macro_inst|controller|serial|shift_data [27];
//wire	\macro_inst|controller|serial|shift_data [28];
//wire	\macro_inst|controller|serial|shift_data [29];
//wire	\macro_inst|controller|serial|shift_data [2];
//wire	\macro_inst|controller|serial|shift_data [30];
//wire	\macro_inst|controller|serial|shift_data [31];
//wire	\macro_inst|controller|serial|shift_data [32];
//wire	\macro_inst|controller|serial|shift_data [33];
//wire	\macro_inst|controller|serial|shift_data [34];
//wire	\macro_inst|controller|serial|shift_data [35];
//wire	\macro_inst|controller|serial|shift_data [36];
//wire	\macro_inst|controller|serial|shift_data [37];
//wire	\macro_inst|controller|serial|shift_data [38];
//wire	\macro_inst|controller|serial|shift_data [39];
//wire	\macro_inst|controller|serial|shift_data [3];
//wire	\macro_inst|controller|serial|shift_data [40];
//wire	\macro_inst|controller|serial|shift_data [41];
//wire	\macro_inst|controller|serial|shift_data [42];
//wire	\macro_inst|controller|serial|shift_data [43];
//wire	\macro_inst|controller|serial|shift_data [44];
//wire	\macro_inst|controller|serial|shift_data [45];
//wire	\macro_inst|controller|serial|shift_data [46];
//wire	\macro_inst|controller|serial|shift_data [47];
wire	\macro_inst|controller|serial|shift_data[47]~1_combout ;
//wire	\macro_inst|controller|serial|shift_data [48];
//wire	\macro_inst|controller|serial|shift_data [49];
//wire	\macro_inst|controller|serial|shift_data [4];
//wire	\macro_inst|controller|serial|shift_data [50];
//wire	\macro_inst|controller|serial|shift_data [51];
//wire	\macro_inst|controller|serial|shift_data [52];
//wire	\macro_inst|controller|serial|shift_data [53];
//wire	\macro_inst|controller|serial|shift_data [54];
//wire	\macro_inst|controller|serial|shift_data [55];
//wire	\macro_inst|controller|serial|shift_data [56];
//wire	\macro_inst|controller|serial|shift_data [57];
//wire	\macro_inst|controller|serial|shift_data [58];
//wire	\macro_inst|controller|serial|shift_data [59];
//wire	\macro_inst|controller|serial|shift_data [5];
//wire	\macro_inst|controller|serial|shift_data [60];
//wire	\macro_inst|controller|serial|shift_data [61];
//wire	\macro_inst|controller|serial|shift_data [62];
//wire	\macro_inst|controller|serial|shift_data [63];
//wire	\macro_inst|controller|serial|shift_data [64];
//wire	\macro_inst|controller|serial|shift_data [65];
//wire	\macro_inst|controller|serial|shift_data [66];
//wire	\macro_inst|controller|serial|shift_data [67];
//wire	\macro_inst|controller|serial|shift_data [68];
//wire	\macro_inst|controller|serial|shift_data [69];
//wire	\macro_inst|controller|serial|shift_data [6];
//wire	\macro_inst|controller|serial|shift_data [70];
//wire	\macro_inst|controller|serial|shift_data [71];
//wire	\macro_inst|controller|serial|shift_data [72];
//wire	\macro_inst|controller|serial|shift_data [73];
//wire	\macro_inst|controller|serial|shift_data [74];
//wire	\macro_inst|controller|serial|shift_data [75];
//wire	\macro_inst|controller|serial|shift_data [76];
//wire	\macro_inst|controller|serial|shift_data [77];
//wire	\macro_inst|controller|serial|shift_data [78];
//wire	\macro_inst|controller|serial|shift_data [79];
//wire	\macro_inst|controller|serial|shift_data [7];
//wire	\macro_inst|controller|serial|shift_data [80];
//wire	\macro_inst|controller|serial|shift_data [81];
//wire	\macro_inst|controller|serial|shift_data [82];
//wire	\macro_inst|controller|serial|shift_data [83];
//wire	\macro_inst|controller|serial|shift_data [84];
//wire	\macro_inst|controller|serial|shift_data [85];
//wire	\macro_inst|controller|serial|shift_data [86];
//wire	\macro_inst|controller|serial|shift_data [87];
//wire	\macro_inst|controller|serial|shift_data [88];
//wire	\macro_inst|controller|serial|shift_data [89];
//wire	\macro_inst|controller|serial|shift_data [8];
//wire	\macro_inst|controller|serial|shift_data [90];
//wire	\macro_inst|controller|serial|shift_data [91];
//wire	\macro_inst|controller|serial|shift_data [92];
//wire	\macro_inst|controller|serial|shift_data [93];
//wire	\macro_inst|controller|serial|shift_data [94];
//wire	\macro_inst|controller|serial|shift_data [95];
//wire	\macro_inst|controller|serial|shift_data [96];
//wire	\macro_inst|controller|serial|shift_data [97];
//wire	\macro_inst|controller|serial|shift_data [98];
//wire	\macro_inst|controller|serial|shift_data [99];
//wire	\macro_inst|controller|serial|shift_data [9];
wire	\macro_inst|controller|serial|shift_data~0_combout ;
wire	\macro_inst|controller|serial|shift_data~100_combout ;
wire	\macro_inst|controller|serial|shift_data~101_combout ;
wire	\macro_inst|controller|serial|shift_data~102_combout ;
wire	\macro_inst|controller|serial|shift_data~103_combout ;
wire	\macro_inst|controller|serial|shift_data~104_combout ;
wire	\macro_inst|controller|serial|shift_data~105_combout ;
wire	\macro_inst|controller|serial|shift_data~106_combout ;
wire	\macro_inst|controller|serial|shift_data~107_combout ;
wire	\macro_inst|controller|serial|shift_data~108_combout ;
wire	\macro_inst|controller|serial|shift_data~109_combout ;
wire	\macro_inst|controller|serial|shift_data~10_combout ;
wire	\macro_inst|controller|serial|shift_data~110_combout ;
wire	\macro_inst|controller|serial|shift_data~111_combout ;
wire	\macro_inst|controller|serial|shift_data~112_combout ;
wire	\macro_inst|controller|serial|shift_data~113_combout ;
wire	\macro_inst|controller|serial|shift_data~114_combout ;
wire	\macro_inst|controller|serial|shift_data~115_combout ;
wire	\macro_inst|controller|serial|shift_data~116_combout ;
wire	\macro_inst|controller|serial|shift_data~117_combout ;
wire	\macro_inst|controller|serial|shift_data~118_combout ;
wire	\macro_inst|controller|serial|shift_data~119_combout ;
wire	\macro_inst|controller|serial|shift_data~11_combout ;
wire	\macro_inst|controller|serial|shift_data~120_combout ;
wire	\macro_inst|controller|serial|shift_data~121_combout ;
wire	\macro_inst|controller|serial|shift_data~122_combout ;
wire	\macro_inst|controller|serial|shift_data~123_combout ;
wire	\macro_inst|controller|serial|shift_data~124_combout ;
wire	\macro_inst|controller|serial|shift_data~125_combout ;
wire	\macro_inst|controller|serial|shift_data~126_combout ;
wire	\macro_inst|controller|serial|shift_data~127_combout ;
wire	\macro_inst|controller|serial|shift_data~128_combout ;
wire	\macro_inst|controller|serial|shift_data~129_combout ;
wire	\macro_inst|controller|serial|shift_data~12_combout ;
wire	\macro_inst|controller|serial|shift_data~130_combout ;
wire	\macro_inst|controller|serial|shift_data~131_combout ;
wire	\macro_inst|controller|serial|shift_data~132_combout ;
wire	\macro_inst|controller|serial|shift_data~133_combout ;
wire	\macro_inst|controller|serial|shift_data~134_combout ;
wire	\macro_inst|controller|serial|shift_data~135_combout ;
wire	\macro_inst|controller|serial|shift_data~136_combout ;
wire	\macro_inst|controller|serial|shift_data~137_combout ;
wire	\macro_inst|controller|serial|shift_data~138_combout ;
wire	\macro_inst|controller|serial|shift_data~139_combout ;
wire	\macro_inst|controller|serial|shift_data~13_combout ;
wire	\macro_inst|controller|serial|shift_data~140_combout ;
wire	\macro_inst|controller|serial|shift_data~141_combout ;
wire	\macro_inst|controller|serial|shift_data~142_combout ;
wire	\macro_inst|controller|serial|shift_data~143_combout ;
wire	\macro_inst|controller|serial|shift_data~144_combout ;
wire	\macro_inst|controller|serial|shift_data~145_combout ;
wire	\macro_inst|controller|serial|shift_data~146_combout ;
wire	\macro_inst|controller|serial|shift_data~147_combout ;
wire	\macro_inst|controller|serial|shift_data~148_combout ;
wire	\macro_inst|controller|serial|shift_data~149_combout ;
wire	\macro_inst|controller|serial|shift_data~14_combout ;
wire	\macro_inst|controller|serial|shift_data~150_combout ;
wire	\macro_inst|controller|serial|shift_data~151_combout ;
wire	\macro_inst|controller|serial|shift_data~152_combout ;
wire	\macro_inst|controller|serial|shift_data~153_combout ;
wire	\macro_inst|controller|serial|shift_data~154_combout ;
wire	\macro_inst|controller|serial|shift_data~155_combout ;
wire	\macro_inst|controller|serial|shift_data~156_combout ;
wire	\macro_inst|controller|serial|shift_data~157_combout ;
wire	\macro_inst|controller|serial|shift_data~158_combout ;
wire	\macro_inst|controller|serial|shift_data~159_combout ;
wire	\macro_inst|controller|serial|shift_data~15_combout ;
wire	\macro_inst|controller|serial|shift_data~160_combout ;
wire	\macro_inst|controller|serial|shift_data~161_combout ;
wire	\macro_inst|controller|serial|shift_data~162_combout ;
wire	\macro_inst|controller|serial|shift_data~163_combout ;
wire	\macro_inst|controller|serial|shift_data~164_combout ;
wire	\macro_inst|controller|serial|shift_data~165_combout ;
wire	\macro_inst|controller|serial|shift_data~166_combout ;
wire	\macro_inst|controller|serial|shift_data~167_combout ;
wire	\macro_inst|controller|serial|shift_data~168_combout ;
wire	\macro_inst|controller|serial|shift_data~169_combout ;
wire	\macro_inst|controller|serial|shift_data~16_combout ;
wire	\macro_inst|controller|serial|shift_data~170_combout ;
wire	\macro_inst|controller|serial|shift_data~171_combout ;
wire	\macro_inst|controller|serial|shift_data~172_combout ;
wire	\macro_inst|controller|serial|shift_data~173_combout ;
wire	\macro_inst|controller|serial|shift_data~174_combout ;
wire	\macro_inst|controller|serial|shift_data~175_combout ;
wire	\macro_inst|controller|serial|shift_data~176_combout ;
wire	\macro_inst|controller|serial|shift_data~177_combout ;
wire	\macro_inst|controller|serial|shift_data~178_combout ;
wire	\macro_inst|controller|serial|shift_data~179_combout ;
wire	\macro_inst|controller|serial|shift_data~17_combout ;
wire	\macro_inst|controller|serial|shift_data~180_combout ;
wire	\macro_inst|controller|serial|shift_data~181_combout ;
wire	\macro_inst|controller|serial|shift_data~182_combout ;
wire	\macro_inst|controller|serial|shift_data~183_combout ;
wire	\macro_inst|controller|serial|shift_data~184_combout ;
wire	\macro_inst|controller|serial|shift_data~185_combout ;
wire	\macro_inst|controller|serial|shift_data~186_combout ;
wire	\macro_inst|controller|serial|shift_data~187_combout ;
wire	\macro_inst|controller|serial|shift_data~188_combout ;
wire	\macro_inst|controller|serial|shift_data~189_combout ;
wire	\macro_inst|controller|serial|shift_data~18_combout ;
wire	\macro_inst|controller|serial|shift_data~190_combout ;
wire	\macro_inst|controller|serial|shift_data~191_combout ;
wire	\macro_inst|controller|serial|shift_data~192_combout ;
wire	\macro_inst|controller|serial|shift_data~19_combout ;
wire	\macro_inst|controller|serial|shift_data~20_combout ;
wire	\macro_inst|controller|serial|shift_data~21_combout ;
wire	\macro_inst|controller|serial|shift_data~22_combout ;
wire	\macro_inst|controller|serial|shift_data~23_combout ;
wire	\macro_inst|controller|serial|shift_data~24_combout ;
wire	\macro_inst|controller|serial|shift_data~25_combout ;
wire	\macro_inst|controller|serial|shift_data~26_combout ;
wire	\macro_inst|controller|serial|shift_data~27_combout ;
wire	\macro_inst|controller|serial|shift_data~28_combout ;
wire	\macro_inst|controller|serial|shift_data~29_combout ;
wire	\macro_inst|controller|serial|shift_data~2_combout ;
wire	\macro_inst|controller|serial|shift_data~30_combout ;
wire	\macro_inst|controller|serial|shift_data~31_combout ;
wire	\macro_inst|controller|serial|shift_data~32_combout ;
wire	\macro_inst|controller|serial|shift_data~33_combout ;
wire	\macro_inst|controller|serial|shift_data~34_combout ;
wire	\macro_inst|controller|serial|shift_data~35_combout ;
wire	\macro_inst|controller|serial|shift_data~36_combout ;
wire	\macro_inst|controller|serial|shift_data~37_combout ;
wire	\macro_inst|controller|serial|shift_data~38_combout ;
wire	\macro_inst|controller|serial|shift_data~39_combout ;
wire	\macro_inst|controller|serial|shift_data~3_combout ;
wire	\macro_inst|controller|serial|shift_data~40_combout ;
wire	\macro_inst|controller|serial|shift_data~41_combout ;
wire	\macro_inst|controller|serial|shift_data~42_combout ;
wire	\macro_inst|controller|serial|shift_data~43_combout ;
wire	\macro_inst|controller|serial|shift_data~44_combout ;
wire	\macro_inst|controller|serial|shift_data~45_combout ;
wire	\macro_inst|controller|serial|shift_data~46_combout ;
wire	\macro_inst|controller|serial|shift_data~47_combout ;
wire	\macro_inst|controller|serial|shift_data~48_combout ;
wire	\macro_inst|controller|serial|shift_data~49_combout ;
wire	\macro_inst|controller|serial|shift_data~4_combout ;
wire	\macro_inst|controller|serial|shift_data~50_combout ;
wire	\macro_inst|controller|serial|shift_data~51_combout ;
wire	\macro_inst|controller|serial|shift_data~52_combout ;
wire	\macro_inst|controller|serial|shift_data~53_combout ;
wire	\macro_inst|controller|serial|shift_data~54_combout ;
wire	\macro_inst|controller|serial|shift_data~55_combout ;
wire	\macro_inst|controller|serial|shift_data~56_combout ;
wire	\macro_inst|controller|serial|shift_data~57_combout ;
wire	\macro_inst|controller|serial|shift_data~58_combout ;
wire	\macro_inst|controller|serial|shift_data~59_combout ;
wire	\macro_inst|controller|serial|shift_data~5_combout ;
wire	\macro_inst|controller|serial|shift_data~60_combout ;
wire	\macro_inst|controller|serial|shift_data~61_combout ;
wire	\macro_inst|controller|serial|shift_data~62_combout ;
wire	\macro_inst|controller|serial|shift_data~63_combout ;
wire	\macro_inst|controller|serial|shift_data~64_combout ;
wire	\macro_inst|controller|serial|shift_data~65_combout ;
wire	\macro_inst|controller|serial|shift_data~66_combout ;
wire	\macro_inst|controller|serial|shift_data~67_combout ;
wire	\macro_inst|controller|serial|shift_data~68_combout ;
wire	\macro_inst|controller|serial|shift_data~69_combout ;
wire	\macro_inst|controller|serial|shift_data~6_combout ;
wire	\macro_inst|controller|serial|shift_data~70_combout ;
wire	\macro_inst|controller|serial|shift_data~71_combout ;
wire	\macro_inst|controller|serial|shift_data~72_combout ;
wire	\macro_inst|controller|serial|shift_data~73_combout ;
wire	\macro_inst|controller|serial|shift_data~74_combout ;
wire	\macro_inst|controller|serial|shift_data~75_combout ;
wire	\macro_inst|controller|serial|shift_data~76_combout ;
wire	\macro_inst|controller|serial|shift_data~77_combout ;
wire	\macro_inst|controller|serial|shift_data~78_combout ;
wire	\macro_inst|controller|serial|shift_data~79_combout ;
wire	\macro_inst|controller|serial|shift_data~7_combout ;
wire	\macro_inst|controller|serial|shift_data~80_combout ;
wire	\macro_inst|controller|serial|shift_data~81_combout ;
wire	\macro_inst|controller|serial|shift_data~82_combout ;
wire	\macro_inst|controller|serial|shift_data~83_combout ;
wire	\macro_inst|controller|serial|shift_data~84_combout ;
wire	\macro_inst|controller|serial|shift_data~85_combout ;
wire	\macro_inst|controller|serial|shift_data~86_combout ;
wire	\macro_inst|controller|serial|shift_data~87_combout ;
wire	\macro_inst|controller|serial|shift_data~88_combout ;
wire	\macro_inst|controller|serial|shift_data~89_combout ;
wire	\macro_inst|controller|serial|shift_data~8_combout ;
wire	\macro_inst|controller|serial|shift_data~90_combout ;
wire	\macro_inst|controller|serial|shift_data~91_combout ;
wire	\macro_inst|controller|serial|shift_data~92_combout ;
wire	\macro_inst|controller|serial|shift_data~93_combout ;
wire	\macro_inst|controller|serial|shift_data~94_combout ;
wire	\macro_inst|controller|serial|shift_data~95_combout ;
wire	\macro_inst|controller|serial|shift_data~96_combout ;
wire	\macro_inst|controller|serial|shift_data~97_combout ;
wire	\macro_inst|controller|serial|shift_data~98_combout ;
wire	\macro_inst|controller|serial|shift_data~99_combout ;
wire	\macro_inst|controller|serial|shift_data~9_combout ;
wire	\macro_inst|controller|serial|shi~0_combout ;
wire	\macro_inst|controller|serial|shi~1_combout ;
wire	\macro_inst|controller|serial|shi~q ;
wire	\macro_inst|controller|serial|state.IDLE~q ;
wire	\macro_inst|controller|serial|state.IDLE~q__SyncLoad_X50_Y1_INV ;
wire	\macro_inst|controller|serial|state.IDLE~q__SyncReset_X51_Y2_INV ;
wire	\macro_inst|controller|serial|state.LATCH~q ;
wire	\macro_inst|controller|serial|state.LOAD~0_combout ;
wire	\macro_inst|controller|serial|state.LOAD~q ;
wire	\macro_inst|controller|serial|state.SHIFT~feeder_combout ;
wire	\macro_inst|controller|serial|state.SHIFT~q ;
wire	\macro_inst|controller|serial|state~14_combout ;
wire	\macro_inst|controller|serial|state~15_combout ;
wire	\macro_inst|controller|serial|sto~0_combout ;
wire	\macro_inst|controller|serial|sto~1_combout ;
wire	\macro_inst|controller|serial|sto~q ;
wire	\macro_inst|controller|sm_pwm|Add0~0_combout ;
wire	\macro_inst|controller|sm_pwm|Add0~1 ;
wire	\macro_inst|controller|sm_pwm|Add0~10_combout ;
wire	\macro_inst|controller|sm_pwm|Add0~11 ;
wire	\macro_inst|controller|sm_pwm|Add0~12_combout ;
wire	\macro_inst|controller|sm_pwm|Add0~13 ;
wire	\macro_inst|controller|sm_pwm|Add0~14_combout ;
wire	\macro_inst|controller|sm_pwm|Add0~2_combout ;
wire	\macro_inst|controller|sm_pwm|Add0~3 ;
wire	\macro_inst|controller|sm_pwm|Add0~4_combout ;
wire	\macro_inst|controller|sm_pwm|Add0~5 ;
wire	\macro_inst|controller|sm_pwm|Add0~6_combout ;
wire	\macro_inst|controller|sm_pwm|Add0~7 ;
wire	\macro_inst|controller|sm_pwm|Add0~8_combout ;
wire	\macro_inst|controller|sm_pwm|Add0~9 ;
wire	\macro_inst|controller|sm_pwm|Decoder0~10_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~11_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~12_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~13_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~14_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~15_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~16_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~17_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~18_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~19_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~20_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~21_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~22_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~23_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~24_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~25_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~26_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~27_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~28_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~29_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~30_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~31_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~32_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~33_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~34_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~35_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~36_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~37_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~38_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~39_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~40_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~41_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~42_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~43_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~44_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~45_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~46_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~47_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~48_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~49_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~4_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~50_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~51_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~52_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~53_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~54_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~55_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~56_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~57_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~58_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~59_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~5_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~60_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~61_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~62_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~63_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~64_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~65_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~66_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~67_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~68_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~69_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~6_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~70_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~71_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~72_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~73_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~74_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~75_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~76_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~77_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~78_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~79_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~7_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~80_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~81_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~8_combout ;
wire	\macro_inst|controller|sm_pwm|Decoder0~9_combout ;
wire	\macro_inst|controller|sm_pwm|Equal0~0_combout ;
wire	\macro_inst|controller|sm_pwm|Equal0~1_combout ;
wire	\macro_inst|controller|sm_pwm|Equal1~0_combout ;
wire	\macro_inst|controller|sm_pwm|Equal1~1_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan0~0_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan10~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan10~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan10~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan10~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan10~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan10~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan10~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan11~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan11~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan11~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan11~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan11~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan11~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan11~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan12~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan12~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan12~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan12~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan12~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan12~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan12~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan13~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan13~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan13~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan13~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan13~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan13~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan13~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan14~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan14~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan14~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan14~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan14~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan14~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan14~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan15~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan15~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan15~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan15~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan15~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan15~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan15~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan16~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan16~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan16~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan16~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan16~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan16~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan16~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan17~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan17~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan17~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan17~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan17~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan17~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan17~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan18~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan18~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan18~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan18~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan18~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan18~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan18~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan19~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan19~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan19~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan19~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan19~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan19~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan19~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan1~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan1~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan1~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan1~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan1~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan1~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan1~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan20~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan20~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan20~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan20~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan20~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan20~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan20~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan21~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan21~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan21~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan21~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan21~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan21~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan21~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan22~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan22~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan22~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan22~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan22~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan22~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan22~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan23~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan23~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan23~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan23~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan23~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan23~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan23~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan24~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan24~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan24~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan24~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan24~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan24~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan24~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan25~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan25~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan25~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan25~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan25~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan25~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan25~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan26~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan26~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan26~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan26~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan26~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan26~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan26~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan27~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan27~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan27~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan27~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan27~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan27~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan27~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan28~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan28~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan28~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan28~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan28~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan28~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan28~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan29~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan29~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan29~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan29~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan29~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan29~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan29~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan2~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan2~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan2~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan2~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan2~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan2~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan2~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan30~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan30~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan30~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan30~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan30~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan30~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan30~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan31~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan31~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan31~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan31~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan31~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan31~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan31~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan32~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan32~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan32~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan32~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan32~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan32~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan32~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan33~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan33~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan33~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan33~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan33~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan33~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan33~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan34~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan34~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan34~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan34~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan34~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan34~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan34~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan35~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan35~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan35~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan35~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan35~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan35~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan35~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan36~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan36~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan36~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan36~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan36~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan36~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan36~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan37~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan37~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan37~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan37~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan37~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan37~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan37~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan38~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan38~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan38~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan38~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan38~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan38~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan38~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan39~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan39~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan39~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan39~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan39~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan39~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan39~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan3~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan3~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan3~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan3~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan3~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan3~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan3~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan40~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan40~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan40~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan40~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan40~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan40~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan40~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan41~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan41~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan41~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan41~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan41~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan41~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan41~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan42~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan42~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan42~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan42~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan42~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan42~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan42~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan43~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan43~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan43~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan43~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan43~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan43~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan43~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan44~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan44~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan44~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan44~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan44~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan44~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan44~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan45~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan45~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan45~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan45~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan45~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan45~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan45~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan46~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan46~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan46~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan46~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan46~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan46~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan46~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan47~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan47~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan47~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan47~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan47~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan47~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan47~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan48~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan48~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan48~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan48~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan48~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan48~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan48~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan49~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan49~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan49~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan49~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan49~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan49~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan49~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan4~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan4~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan4~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan4~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan4~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan4~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan4~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan50~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan50~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan50~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan50~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan50~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan50~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan50~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan51~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan51~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan51~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan51~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan51~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan51~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan51~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan52~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan52~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan52~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan52~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan52~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan52~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan52~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan53~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan53~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan53~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan53~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan53~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan53~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan53~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan54~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan54~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan54~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan54~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan54~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan54~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan54~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan55~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan55~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan55~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan55~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan55~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan55~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan55~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan56~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan56~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan56~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan56~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan56~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan56~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan56~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan57~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan57~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan57~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan57~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan57~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan57~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan57~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan58~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan58~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan58~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan58~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan58~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan58~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan58~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan59~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan59~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan59~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan59~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan59~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan59~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan59~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan5~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan5~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan5~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan5~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan5~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan5~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan5~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan60~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan60~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan60~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan60~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan60~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan60~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan60~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan61~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan61~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan61~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan61~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan61~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan61~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan61~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan62~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan62~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan62~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan62~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan62~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan62~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan62~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan63~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan63~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan63~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan63~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan63~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan63~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan63~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan64~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan64~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan64~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan64~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan64~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan64~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan64~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan65~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan65~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan65~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan65~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan65~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan65~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan65~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan66~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan66~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan66~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan66~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan66~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan66~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan66~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan67~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan67~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan67~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan67~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan67~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan67~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan67~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan68~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan68~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan68~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan68~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan68~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan68~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan68~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan69~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan69~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan69~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan69~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan69~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan69~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan69~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan6~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan6~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan6~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan6~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan6~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan6~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan6~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan70~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan70~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan70~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan70~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan70~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan70~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan70~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan71~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan71~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan71~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan71~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan71~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan71~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan71~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan72~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan72~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan72~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan72~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan72~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan72~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan72~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan73~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan73~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan73~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan73~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan73~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan73~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan73~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan74~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan74~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan74~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan74~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan74~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan74~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan74~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan75~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan75~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan75~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan75~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan75~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan75~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan75~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan76~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan76~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan76~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan76~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan76~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan76~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan76~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan77~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan77~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan77~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan77~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan77~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan77~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan77~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan78~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan78~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan78~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan78~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan78~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan78~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan78~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan79~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan79~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan79~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan79~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan79~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan79~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan79~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan7~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan7~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan7~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan7~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan7~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan7~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan7~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan80~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan80~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan80~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan80~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan80~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan80~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan80~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan81~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan81~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan81~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan81~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan81~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan81~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan81~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan82~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan82~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan82~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan82~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan82~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan82~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan82~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan83~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan83~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan83~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan83~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan83~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan83~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan83~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan84~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan84~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan84~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan84~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan84~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan84~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan84~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan85~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan85~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan85~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan85~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan85~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan85~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan85~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan86~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan86~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan86~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan86~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan86~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan86~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan86~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan87~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan87~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan87~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan87~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan87~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan87~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan87~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan88~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan88~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan88~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan88~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan88~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan88~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan88~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan89~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan89~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan89~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan89~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan89~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan89~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan89~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan8~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan8~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan8~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan8~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan8~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan8~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan8~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan90~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan90~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan90~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan90~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan90~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan90~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan90~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan91~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan91~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan91~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan91~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan91~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan91~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan91~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan92~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan92~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan92~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan92~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan92~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan92~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan92~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan93~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan93~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan93~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan93~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan93~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan93~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan93~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan94~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan94~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan94~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan94~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan94~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan94~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan94~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan95~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan95~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan95~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan95~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan95~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan95~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan95~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan96~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan96~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan96~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan96~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan96~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan96~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan96~9_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan9~11_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan9~12_combout ;
wire	\macro_inst|controller|sm_pwm|LessThan9~1_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan9~3_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan9~5_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan9~7_cout ;
wire	\macro_inst|controller|sm_pwm|LessThan9~9_cout ;
wire	[191:0] \macro_inst|controller|sm_pwm|data ;
//wire	\macro_inst|controller|sm_pwm|data [0];
//wire	\macro_inst|controller|sm_pwm|data [100];
//wire	\macro_inst|controller|sm_pwm|data [101];
//wire	\macro_inst|controller|sm_pwm|data [102];
//wire	\macro_inst|controller|sm_pwm|data [103];
//wire	\macro_inst|controller|sm_pwm|data [104];
//wire	\macro_inst|controller|sm_pwm|data [105];
//wire	\macro_inst|controller|sm_pwm|data [106];
//wire	\macro_inst|controller|sm_pwm|data [107];
//wire	\macro_inst|controller|sm_pwm|data [108];
//wire	\macro_inst|controller|sm_pwm|data [109];
//wire	\macro_inst|controller|sm_pwm|data [10];
//wire	\macro_inst|controller|sm_pwm|data [110];
//wire	\macro_inst|controller|sm_pwm|data [111];
//wire	\macro_inst|controller|sm_pwm|data [112];
//wire	\macro_inst|controller|sm_pwm|data [113];
//wire	\macro_inst|controller|sm_pwm|data [114];
//wire	\macro_inst|controller|sm_pwm|data [115];
//wire	\macro_inst|controller|sm_pwm|data [116];
//wire	\macro_inst|controller|sm_pwm|data [117];
//wire	\macro_inst|controller|sm_pwm|data [118];
//wire	\macro_inst|controller|sm_pwm|data [119];
//wire	\macro_inst|controller|sm_pwm|data [11];
//wire	\macro_inst|controller|sm_pwm|data [120];
//wire	\macro_inst|controller|sm_pwm|data [121];
//wire	\macro_inst|controller|sm_pwm|data [122];
//wire	\macro_inst|controller|sm_pwm|data [123];
//wire	\macro_inst|controller|sm_pwm|data [124];
//wire	\macro_inst|controller|sm_pwm|data [125];
//wire	\macro_inst|controller|sm_pwm|data [126];
//wire	\macro_inst|controller|sm_pwm|data [127];
//wire	\macro_inst|controller|sm_pwm|data [128];
//wire	\macro_inst|controller|sm_pwm|data [129];
//wire	\macro_inst|controller|sm_pwm|data [12];
//wire	\macro_inst|controller|sm_pwm|data [130];
//wire	\macro_inst|controller|sm_pwm|data [131];
//wire	\macro_inst|controller|sm_pwm|data [132];
//wire	\macro_inst|controller|sm_pwm|data [133];
//wire	\macro_inst|controller|sm_pwm|data [134];
//wire	\macro_inst|controller|sm_pwm|data [135];
//wire	\macro_inst|controller|sm_pwm|data [136];
//wire	\macro_inst|controller|sm_pwm|data [137];
//wire	\macro_inst|controller|sm_pwm|data [138];
//wire	\macro_inst|controller|sm_pwm|data [139];
//wire	\macro_inst|controller|sm_pwm|data [13];
//wire	\macro_inst|controller|sm_pwm|data [140];
//wire	\macro_inst|controller|sm_pwm|data [141];
//wire	\macro_inst|controller|sm_pwm|data [142];
//wire	\macro_inst|controller|sm_pwm|data [143];
//wire	\macro_inst|controller|sm_pwm|data [144];
//wire	\macro_inst|controller|sm_pwm|data [145];
//wire	\macro_inst|controller|sm_pwm|data [146];
//wire	\macro_inst|controller|sm_pwm|data [147];
//wire	\macro_inst|controller|sm_pwm|data [148];
//wire	\macro_inst|controller|sm_pwm|data [149];
//wire	\macro_inst|controller|sm_pwm|data [14];
//wire	\macro_inst|controller|sm_pwm|data [150];
//wire	\macro_inst|controller|sm_pwm|data [151];
//wire	\macro_inst|controller|sm_pwm|data [152];
//wire	\macro_inst|controller|sm_pwm|data [153];
//wire	\macro_inst|controller|sm_pwm|data [154];
//wire	\macro_inst|controller|sm_pwm|data [155];
//wire	\macro_inst|controller|sm_pwm|data [156];
//wire	\macro_inst|controller|sm_pwm|data [157];
//wire	\macro_inst|controller|sm_pwm|data [158];
//wire	\macro_inst|controller|sm_pwm|data [159];
//wire	\macro_inst|controller|sm_pwm|data [15];
//wire	\macro_inst|controller|sm_pwm|data [160];
//wire	\macro_inst|controller|sm_pwm|data [161];
//wire	\macro_inst|controller|sm_pwm|data [162];
//wire	\macro_inst|controller|sm_pwm|data [163];
//wire	\macro_inst|controller|sm_pwm|data [164];
//wire	\macro_inst|controller|sm_pwm|data [165];
//wire	\macro_inst|controller|sm_pwm|data [166];
//wire	\macro_inst|controller|sm_pwm|data [167];
//wire	\macro_inst|controller|sm_pwm|data [168];
//wire	\macro_inst|controller|sm_pwm|data [169];
//wire	\macro_inst|controller|sm_pwm|data [16];
//wire	\macro_inst|controller|sm_pwm|data [170];
//wire	\macro_inst|controller|sm_pwm|data [171];
//wire	\macro_inst|controller|sm_pwm|data [172];
//wire	\macro_inst|controller|sm_pwm|data [173];
//wire	\macro_inst|controller|sm_pwm|data [174];
//wire	\macro_inst|controller|sm_pwm|data [175];
//wire	\macro_inst|controller|sm_pwm|data [176];
//wire	\macro_inst|controller|sm_pwm|data [177];
//wire	\macro_inst|controller|sm_pwm|data [178];
//wire	\macro_inst|controller|sm_pwm|data [179];
//wire	\macro_inst|controller|sm_pwm|data [17];
//wire	\macro_inst|controller|sm_pwm|data [180];
//wire	\macro_inst|controller|sm_pwm|data [181];
//wire	\macro_inst|controller|sm_pwm|data [182];
//wire	\macro_inst|controller|sm_pwm|data [183];
//wire	\macro_inst|controller|sm_pwm|data [184];
//wire	\macro_inst|controller|sm_pwm|data [185];
//wire	\macro_inst|controller|sm_pwm|data [186];
//wire	\macro_inst|controller|sm_pwm|data [187];
//wire	\macro_inst|controller|sm_pwm|data [188];
//wire	\macro_inst|controller|sm_pwm|data [189];
//wire	\macro_inst|controller|sm_pwm|data [18];
//wire	\macro_inst|controller|sm_pwm|data [190];
//wire	\macro_inst|controller|sm_pwm|data [191];
//wire	\macro_inst|controller|sm_pwm|data [19];
//wire	\macro_inst|controller|sm_pwm|data [1];
//wire	\macro_inst|controller|sm_pwm|data [20];
//wire	\macro_inst|controller|sm_pwm|data [21];
//wire	\macro_inst|controller|sm_pwm|data [22];
//wire	\macro_inst|controller|sm_pwm|data [23];
//wire	\macro_inst|controller|sm_pwm|data [24];
//wire	\macro_inst|controller|sm_pwm|data [25];
//wire	\macro_inst|controller|sm_pwm|data [26];
//wire	\macro_inst|controller|sm_pwm|data [27];
//wire	\macro_inst|controller|sm_pwm|data [28];
//wire	\macro_inst|controller|sm_pwm|data [29];
//wire	\macro_inst|controller|sm_pwm|data [2];
//wire	\macro_inst|controller|sm_pwm|data [30];
//wire	\macro_inst|controller|sm_pwm|data [31];
//wire	\macro_inst|controller|sm_pwm|data [32];
//wire	\macro_inst|controller|sm_pwm|data [33];
//wire	\macro_inst|controller|sm_pwm|data [34];
//wire	\macro_inst|controller|sm_pwm|data [35];
//wire	\macro_inst|controller|sm_pwm|data [36];
//wire	\macro_inst|controller|sm_pwm|data [37];
//wire	\macro_inst|controller|sm_pwm|data [38];
//wire	\macro_inst|controller|sm_pwm|data [39];
//wire	\macro_inst|controller|sm_pwm|data [3];
//wire	\macro_inst|controller|sm_pwm|data [40];
//wire	\macro_inst|controller|sm_pwm|data [41];
//wire	\macro_inst|controller|sm_pwm|data [42];
//wire	\macro_inst|controller|sm_pwm|data [43];
//wire	\macro_inst|controller|sm_pwm|data [44];
//wire	\macro_inst|controller|sm_pwm|data [45];
//wire	\macro_inst|controller|sm_pwm|data [46];
//wire	\macro_inst|controller|sm_pwm|data [47];
//wire	\macro_inst|controller|sm_pwm|data [48];
//wire	\macro_inst|controller|sm_pwm|data [49];
//wire	\macro_inst|controller|sm_pwm|data [4];
//wire	\macro_inst|controller|sm_pwm|data [50];
//wire	\macro_inst|controller|sm_pwm|data [51];
//wire	\macro_inst|controller|sm_pwm|data [52];
//wire	\macro_inst|controller|sm_pwm|data [53];
//wire	\macro_inst|controller|sm_pwm|data [54];
//wire	\macro_inst|controller|sm_pwm|data [55];
//wire	\macro_inst|controller|sm_pwm|data [56];
//wire	\macro_inst|controller|sm_pwm|data [57];
//wire	\macro_inst|controller|sm_pwm|data [58];
//wire	\macro_inst|controller|sm_pwm|data [59];
//wire	\macro_inst|controller|sm_pwm|data [5];
//wire	\macro_inst|controller|sm_pwm|data [60];
//wire	\macro_inst|controller|sm_pwm|data [61];
//wire	\macro_inst|controller|sm_pwm|data [62];
//wire	\macro_inst|controller|sm_pwm|data [63];
//wire	\macro_inst|controller|sm_pwm|data [64];
//wire	\macro_inst|controller|sm_pwm|data [65];
//wire	\macro_inst|controller|sm_pwm|data [66];
//wire	\macro_inst|controller|sm_pwm|data [67];
//wire	\macro_inst|controller|sm_pwm|data [68];
//wire	\macro_inst|controller|sm_pwm|data [69];
//wire	\macro_inst|controller|sm_pwm|data [6];
//wire	\macro_inst|controller|sm_pwm|data [70];
//wire	\macro_inst|controller|sm_pwm|data [71];
//wire	\macro_inst|controller|sm_pwm|data [72];
//wire	\macro_inst|controller|sm_pwm|data [73];
//wire	\macro_inst|controller|sm_pwm|data [74];
//wire	\macro_inst|controller|sm_pwm|data [75];
//wire	\macro_inst|controller|sm_pwm|data [76];
//wire	\macro_inst|controller|sm_pwm|data [77];
//wire	\macro_inst|controller|sm_pwm|data [78];
//wire	\macro_inst|controller|sm_pwm|data [79];
//wire	\macro_inst|controller|sm_pwm|data [7];
//wire	\macro_inst|controller|sm_pwm|data [80];
//wire	\macro_inst|controller|sm_pwm|data [81];
//wire	\macro_inst|controller|sm_pwm|data [82];
//wire	\macro_inst|controller|sm_pwm|data [83];
//wire	\macro_inst|controller|sm_pwm|data [84];
//wire	\macro_inst|controller|sm_pwm|data [85];
//wire	\macro_inst|controller|sm_pwm|data [86];
//wire	\macro_inst|controller|sm_pwm|data [87];
//wire	\macro_inst|controller|sm_pwm|data [88];
//wire	\macro_inst|controller|sm_pwm|data [89];
//wire	\macro_inst|controller|sm_pwm|data [8];
//wire	\macro_inst|controller|sm_pwm|data [90];
//wire	\macro_inst|controller|sm_pwm|data [91];
//wire	\macro_inst|controller|sm_pwm|data [92];
//wire	\macro_inst|controller|sm_pwm|data [93];
//wire	\macro_inst|controller|sm_pwm|data [94];
//wire	\macro_inst|controller|sm_pwm|data [95];
//wire	\macro_inst|controller|sm_pwm|data [96];
//wire	\macro_inst|controller|sm_pwm|data [97];
//wire	\macro_inst|controller|sm_pwm|data [98];
//wire	\macro_inst|controller|sm_pwm|data [99];
//wire	\macro_inst|controller|sm_pwm|data [9];
wire	\macro_inst|controller|sm_pwm|data~0_combout ;
wire	\macro_inst|controller|sm_pwm|data~100_combout ;
wire	\macro_inst|controller|sm_pwm|data~101_combout ;
wire	\macro_inst|controller|sm_pwm|data~102_combout ;
wire	\macro_inst|controller|sm_pwm|data~103_combout ;
wire	\macro_inst|controller|sm_pwm|data~104_combout ;
wire	\macro_inst|controller|sm_pwm|data~105_combout ;
wire	\macro_inst|controller|sm_pwm|data~106_combout ;
wire	\macro_inst|controller|sm_pwm|data~107_combout ;
wire	\macro_inst|controller|sm_pwm|data~108_combout ;
wire	\macro_inst|controller|sm_pwm|data~109_combout ;
wire	\macro_inst|controller|sm_pwm|data~10_combout ;
wire	\macro_inst|controller|sm_pwm|data~110_combout ;
wire	\macro_inst|controller|sm_pwm|data~111_combout ;
wire	\macro_inst|controller|sm_pwm|data~112_combout ;
wire	\macro_inst|controller|sm_pwm|data~113_combout ;
wire	\macro_inst|controller|sm_pwm|data~114_combout ;
wire	\macro_inst|controller|sm_pwm|data~115_combout ;
wire	\macro_inst|controller|sm_pwm|data~116_combout ;
wire	\macro_inst|controller|sm_pwm|data~117_combout ;
wire	\macro_inst|controller|sm_pwm|data~118_combout ;
wire	\macro_inst|controller|sm_pwm|data~119_combout ;
wire	\macro_inst|controller|sm_pwm|data~11_combout ;
wire	\macro_inst|controller|sm_pwm|data~120_combout ;
wire	\macro_inst|controller|sm_pwm|data~121_combout ;
wire	\macro_inst|controller|sm_pwm|data~122_combout ;
wire	\macro_inst|controller|sm_pwm|data~123_combout ;
wire	\macro_inst|controller|sm_pwm|data~124_combout ;
wire	\macro_inst|controller|sm_pwm|data~125_combout ;
wire	\macro_inst|controller|sm_pwm|data~126_combout ;
wire	\macro_inst|controller|sm_pwm|data~127_combout ;
wire	\macro_inst|controller|sm_pwm|data~128_combout ;
wire	\macro_inst|controller|sm_pwm|data~129_combout ;
wire	\macro_inst|controller|sm_pwm|data~12_combout ;
wire	\macro_inst|controller|sm_pwm|data~130_combout ;
wire	\macro_inst|controller|sm_pwm|data~131_combout ;
wire	\macro_inst|controller|sm_pwm|data~132_combout ;
wire	\macro_inst|controller|sm_pwm|data~133_combout ;
wire	\macro_inst|controller|sm_pwm|data~134_combout ;
wire	\macro_inst|controller|sm_pwm|data~135_combout ;
wire	\macro_inst|controller|sm_pwm|data~136_combout ;
wire	\macro_inst|controller|sm_pwm|data~137_combout ;
wire	\macro_inst|controller|sm_pwm|data~138_combout ;
wire	\macro_inst|controller|sm_pwm|data~139_combout ;
wire	\macro_inst|controller|sm_pwm|data~13_combout ;
wire	\macro_inst|controller|sm_pwm|data~140_combout ;
wire	\macro_inst|controller|sm_pwm|data~141_combout ;
wire	\macro_inst|controller|sm_pwm|data~142_combout ;
wire	\macro_inst|controller|sm_pwm|data~143_combout ;
wire	\macro_inst|controller|sm_pwm|data~144_combout ;
wire	\macro_inst|controller|sm_pwm|data~145_combout ;
wire	\macro_inst|controller|sm_pwm|data~146_combout ;
wire	\macro_inst|controller|sm_pwm|data~147_combout ;
wire	\macro_inst|controller|sm_pwm|data~148_combout ;
wire	\macro_inst|controller|sm_pwm|data~149_combout ;
wire	\macro_inst|controller|sm_pwm|data~14_combout ;
wire	\macro_inst|controller|sm_pwm|data~150_combout ;
wire	\macro_inst|controller|sm_pwm|data~151_combout ;
wire	\macro_inst|controller|sm_pwm|data~152_combout ;
wire	\macro_inst|controller|sm_pwm|data~153_combout ;
wire	\macro_inst|controller|sm_pwm|data~154_combout ;
wire	\macro_inst|controller|sm_pwm|data~155_combout ;
wire	\macro_inst|controller|sm_pwm|data~156_combout ;
wire	\macro_inst|controller|sm_pwm|data~157_combout ;
wire	\macro_inst|controller|sm_pwm|data~158_combout ;
wire	\macro_inst|controller|sm_pwm|data~159_combout ;
wire	\macro_inst|controller|sm_pwm|data~15_combout ;
wire	\macro_inst|controller|sm_pwm|data~160_combout ;
wire	\macro_inst|controller|sm_pwm|data~161_combout ;
wire	\macro_inst|controller|sm_pwm|data~162_combout ;
wire	\macro_inst|controller|sm_pwm|data~163_combout ;
wire	\macro_inst|controller|sm_pwm|data~164_combout ;
wire	\macro_inst|controller|sm_pwm|data~165_combout ;
wire	\macro_inst|controller|sm_pwm|data~166_combout ;
wire	\macro_inst|controller|sm_pwm|data~167_combout ;
wire	\macro_inst|controller|sm_pwm|data~168_combout ;
wire	\macro_inst|controller|sm_pwm|data~169_combout ;
wire	\macro_inst|controller|sm_pwm|data~16_combout ;
wire	\macro_inst|controller|sm_pwm|data~170_combout ;
wire	\macro_inst|controller|sm_pwm|data~171_combout ;
wire	\macro_inst|controller|sm_pwm|data~172_combout ;
wire	\macro_inst|controller|sm_pwm|data~173_combout ;
wire	\macro_inst|controller|sm_pwm|data~174_combout ;
wire	\macro_inst|controller|sm_pwm|data~175_combout ;
wire	\macro_inst|controller|sm_pwm|data~176_combout ;
wire	\macro_inst|controller|sm_pwm|data~177_combout ;
wire	\macro_inst|controller|sm_pwm|data~178_combout ;
wire	\macro_inst|controller|sm_pwm|data~179_combout ;
wire	\macro_inst|controller|sm_pwm|data~17_combout ;
wire	\macro_inst|controller|sm_pwm|data~180_combout ;
wire	\macro_inst|controller|sm_pwm|data~181_combout ;
wire	\macro_inst|controller|sm_pwm|data~182_combout ;
wire	\macro_inst|controller|sm_pwm|data~183_combout ;
wire	\macro_inst|controller|sm_pwm|data~184_combout ;
wire	\macro_inst|controller|sm_pwm|data~185_combout ;
wire	\macro_inst|controller|sm_pwm|data~186_combout ;
wire	\macro_inst|controller|sm_pwm|data~187_combout ;
wire	\macro_inst|controller|sm_pwm|data~188_combout ;
wire	\macro_inst|controller|sm_pwm|data~189_combout ;
wire	\macro_inst|controller|sm_pwm|data~18_combout ;
wire	\macro_inst|controller|sm_pwm|data~190_combout ;
wire	\macro_inst|controller|sm_pwm|data~191_combout ;
wire	\macro_inst|controller|sm_pwm|data~192_combout ;
wire	\macro_inst|controller|sm_pwm|data~193_combout ;
wire	\macro_inst|controller|sm_pwm|data~194_combout ;
wire	\macro_inst|controller|sm_pwm|data~195_combout ;
wire	\macro_inst|controller|sm_pwm|data~196_combout ;
wire	\macro_inst|controller|sm_pwm|data~197_combout ;
wire	\macro_inst|controller|sm_pwm|data~198_combout ;
wire	\macro_inst|controller|sm_pwm|data~199_combout ;
wire	\macro_inst|controller|sm_pwm|data~19_combout ;
wire	\macro_inst|controller|sm_pwm|data~1_combout ;
wire	\macro_inst|controller|sm_pwm|data~200_combout ;
wire	\macro_inst|controller|sm_pwm|data~201_combout ;
wire	\macro_inst|controller|sm_pwm|data~202_combout ;
wire	\macro_inst|controller|sm_pwm|data~203_combout ;
wire	\macro_inst|controller|sm_pwm|data~204_combout ;
wire	\macro_inst|controller|sm_pwm|data~205_combout ;
wire	\macro_inst|controller|sm_pwm|data~206_combout ;
wire	\macro_inst|controller|sm_pwm|data~207_combout ;
wire	\macro_inst|controller|sm_pwm|data~208_combout ;
wire	\macro_inst|controller|sm_pwm|data~209_combout ;
wire	\macro_inst|controller|sm_pwm|data~20_combout ;
wire	\macro_inst|controller|sm_pwm|data~210_combout ;
wire	\macro_inst|controller|sm_pwm|data~211_combout ;
wire	\macro_inst|controller|sm_pwm|data~212_combout ;
wire	\macro_inst|controller|sm_pwm|data~213_combout ;
wire	\macro_inst|controller|sm_pwm|data~214_combout ;
wire	\macro_inst|controller|sm_pwm|data~215_combout ;
wire	\macro_inst|controller|sm_pwm|data~216_combout ;
wire	\macro_inst|controller|sm_pwm|data~217_combout ;
wire	\macro_inst|controller|sm_pwm|data~218_combout ;
wire	\macro_inst|controller|sm_pwm|data~219_combout ;
wire	\macro_inst|controller|sm_pwm|data~21_combout ;
wire	\macro_inst|controller|sm_pwm|data~220_combout ;
wire	\macro_inst|controller|sm_pwm|data~221_combout ;
wire	\macro_inst|controller|sm_pwm|data~222_combout ;
wire	\macro_inst|controller|sm_pwm|data~223_combout ;
wire	\macro_inst|controller|sm_pwm|data~224_combout ;
wire	\macro_inst|controller|sm_pwm|data~225_combout ;
wire	\macro_inst|controller|sm_pwm|data~226_combout ;
wire	\macro_inst|controller|sm_pwm|data~227_combout ;
wire	\macro_inst|controller|sm_pwm|data~228_combout ;
wire	\macro_inst|controller|sm_pwm|data~229_combout ;
wire	\macro_inst|controller|sm_pwm|data~22_combout ;
wire	\macro_inst|controller|sm_pwm|data~230_combout ;
wire	\macro_inst|controller|sm_pwm|data~231_combout ;
wire	\macro_inst|controller|sm_pwm|data~232_combout ;
wire	\macro_inst|controller|sm_pwm|data~233_combout ;
wire	\macro_inst|controller|sm_pwm|data~234_combout ;
wire	\macro_inst|controller|sm_pwm|data~235_combout ;
wire	\macro_inst|controller|sm_pwm|data~236_combout ;
wire	\macro_inst|controller|sm_pwm|data~237_combout ;
wire	\macro_inst|controller|sm_pwm|data~238_combout ;
wire	\macro_inst|controller|sm_pwm|data~239_combout ;
wire	\macro_inst|controller|sm_pwm|data~23_combout ;
wire	\macro_inst|controller|sm_pwm|data~240_combout ;
wire	\macro_inst|controller|sm_pwm|data~241_combout ;
wire	\macro_inst|controller|sm_pwm|data~242_combout ;
wire	\macro_inst|controller|sm_pwm|data~243_combout ;
wire	\macro_inst|controller|sm_pwm|data~244_combout ;
wire	\macro_inst|controller|sm_pwm|data~245_combout ;
wire	\macro_inst|controller|sm_pwm|data~246_combout ;
wire	\macro_inst|controller|sm_pwm|data~247_combout ;
wire	\macro_inst|controller|sm_pwm|data~248_combout ;
wire	\macro_inst|controller|sm_pwm|data~249_combout ;
wire	\macro_inst|controller|sm_pwm|data~24_combout ;
wire	\macro_inst|controller|sm_pwm|data~250_combout ;
wire	\macro_inst|controller|sm_pwm|data~251_combout ;
wire	\macro_inst|controller|sm_pwm|data~252_combout ;
wire	\macro_inst|controller|sm_pwm|data~253_combout ;
wire	\macro_inst|controller|sm_pwm|data~254_combout ;
wire	\macro_inst|controller|sm_pwm|data~255_combout ;
wire	\macro_inst|controller|sm_pwm|data~256_combout ;
wire	\macro_inst|controller|sm_pwm|data~257_combout ;
wire	\macro_inst|controller|sm_pwm|data~258_combout ;
wire	\macro_inst|controller|sm_pwm|data~259_combout ;
wire	\macro_inst|controller|sm_pwm|data~25_combout ;
wire	\macro_inst|controller|sm_pwm|data~260_combout ;
wire	\macro_inst|controller|sm_pwm|data~261_combout ;
wire	\macro_inst|controller|sm_pwm|data~262_combout ;
wire	\macro_inst|controller|sm_pwm|data~263_combout ;
wire	\macro_inst|controller|sm_pwm|data~264_combout ;
wire	\macro_inst|controller|sm_pwm|data~265_combout ;
wire	\macro_inst|controller|sm_pwm|data~266_combout ;
wire	\macro_inst|controller|sm_pwm|data~267_combout ;
wire	\macro_inst|controller|sm_pwm|data~268_combout ;
wire	\macro_inst|controller|sm_pwm|data~269_combout ;
wire	\macro_inst|controller|sm_pwm|data~26_combout ;
wire	\macro_inst|controller|sm_pwm|data~270_combout ;
wire	\macro_inst|controller|sm_pwm|data~271_combout ;
wire	\macro_inst|controller|sm_pwm|data~272_combout ;
wire	\macro_inst|controller|sm_pwm|data~273_combout ;
wire	\macro_inst|controller|sm_pwm|data~274_combout ;
wire	\macro_inst|controller|sm_pwm|data~275_combout ;
wire	\macro_inst|controller|sm_pwm|data~276_combout ;
wire	\macro_inst|controller|sm_pwm|data~277_combout ;
wire	\macro_inst|controller|sm_pwm|data~278_combout ;
wire	\macro_inst|controller|sm_pwm|data~279_combout ;
wire	\macro_inst|controller|sm_pwm|data~27_combout ;
wire	\macro_inst|controller|sm_pwm|data~280_combout ;
wire	\macro_inst|controller|sm_pwm|data~281_combout ;
wire	\macro_inst|controller|sm_pwm|data~282_combout ;
wire	\macro_inst|controller|sm_pwm|data~283_combout ;
wire	\macro_inst|controller|sm_pwm|data~284_combout ;
wire	\macro_inst|controller|sm_pwm|data~285_combout ;
wire	\macro_inst|controller|sm_pwm|data~286_combout ;
wire	\macro_inst|controller|sm_pwm|data~287_combout ;
wire	\macro_inst|controller|sm_pwm|data~28_combout ;
wire	\macro_inst|controller|sm_pwm|data~29_combout ;
wire	\macro_inst|controller|sm_pwm|data~2_combout ;
wire	\macro_inst|controller|sm_pwm|data~30_combout ;
wire	\macro_inst|controller|sm_pwm|data~31_combout ;
wire	\macro_inst|controller|sm_pwm|data~32_combout ;
wire	\macro_inst|controller|sm_pwm|data~33_combout ;
wire	\macro_inst|controller|sm_pwm|data~34_combout ;
wire	\macro_inst|controller|sm_pwm|data~35_combout ;
wire	\macro_inst|controller|sm_pwm|data~36_combout ;
wire	\macro_inst|controller|sm_pwm|data~37_combout ;
wire	\macro_inst|controller|sm_pwm|data~38_combout ;
wire	\macro_inst|controller|sm_pwm|data~39_combout ;
wire	\macro_inst|controller|sm_pwm|data~3_combout ;
wire	\macro_inst|controller|sm_pwm|data~40_combout ;
wire	\macro_inst|controller|sm_pwm|data~41_combout ;
wire	\macro_inst|controller|sm_pwm|data~42_combout ;
wire	\macro_inst|controller|sm_pwm|data~43_combout ;
wire	\macro_inst|controller|sm_pwm|data~44_combout ;
wire	\macro_inst|controller|sm_pwm|data~45_combout ;
wire	\macro_inst|controller|sm_pwm|data~46_combout ;
wire	\macro_inst|controller|sm_pwm|data~47_combout ;
wire	\macro_inst|controller|sm_pwm|data~48_combout ;
wire	\macro_inst|controller|sm_pwm|data~49_combout ;
wire	\macro_inst|controller|sm_pwm|data~4_combout ;
wire	\macro_inst|controller|sm_pwm|data~50_combout ;
wire	\macro_inst|controller|sm_pwm|data~51_combout ;
wire	\macro_inst|controller|sm_pwm|data~52_combout ;
wire	\macro_inst|controller|sm_pwm|data~53_combout ;
wire	\macro_inst|controller|sm_pwm|data~54_combout ;
wire	\macro_inst|controller|sm_pwm|data~55_combout ;
wire	\macro_inst|controller|sm_pwm|data~56_combout ;
wire	\macro_inst|controller|sm_pwm|data~57_combout ;
wire	\macro_inst|controller|sm_pwm|data~58_combout ;
wire	\macro_inst|controller|sm_pwm|data~59_combout ;
wire	\macro_inst|controller|sm_pwm|data~5_combout ;
wire	\macro_inst|controller|sm_pwm|data~60_combout ;
wire	\macro_inst|controller|sm_pwm|data~61_combout ;
wire	\macro_inst|controller|sm_pwm|data~62_combout ;
wire	\macro_inst|controller|sm_pwm|data~63_combout ;
wire	\macro_inst|controller|sm_pwm|data~64_combout ;
wire	\macro_inst|controller|sm_pwm|data~65_combout ;
wire	\macro_inst|controller|sm_pwm|data~66_combout ;
wire	\macro_inst|controller|sm_pwm|data~67_combout ;
wire	\macro_inst|controller|sm_pwm|data~68_combout ;
wire	\macro_inst|controller|sm_pwm|data~69_combout ;
wire	\macro_inst|controller|sm_pwm|data~6_combout ;
wire	\macro_inst|controller|sm_pwm|data~70_combout ;
wire	\macro_inst|controller|sm_pwm|data~71_combout ;
wire	\macro_inst|controller|sm_pwm|data~72_combout ;
wire	\macro_inst|controller|sm_pwm|data~73_combout ;
wire	\macro_inst|controller|sm_pwm|data~74_combout ;
wire	\macro_inst|controller|sm_pwm|data~75_combout ;
wire	\macro_inst|controller|sm_pwm|data~76_combout ;
wire	\macro_inst|controller|sm_pwm|data~77_combout ;
wire	\macro_inst|controller|sm_pwm|data~78_combout ;
wire	\macro_inst|controller|sm_pwm|data~79_combout ;
wire	\macro_inst|controller|sm_pwm|data~7_combout ;
wire	\macro_inst|controller|sm_pwm|data~80_combout ;
wire	\macro_inst|controller|sm_pwm|data~81_combout ;
wire	\macro_inst|controller|sm_pwm|data~82_combout ;
wire	\macro_inst|controller|sm_pwm|data~83_combout ;
wire	\macro_inst|controller|sm_pwm|data~84_combout ;
wire	\macro_inst|controller|sm_pwm|data~85_combout ;
wire	\macro_inst|controller|sm_pwm|data~86_combout ;
wire	\macro_inst|controller|sm_pwm|data~87_combout ;
wire	\macro_inst|controller|sm_pwm|data~88_combout ;
wire	\macro_inst|controller|sm_pwm|data~89_combout ;
wire	\macro_inst|controller|sm_pwm|data~8_combout ;
wire	\macro_inst|controller|sm_pwm|data~90_combout ;
wire	\macro_inst|controller|sm_pwm|data~91_combout ;
wire	\macro_inst|controller|sm_pwm|data~92_combout ;
wire	\macro_inst|controller|sm_pwm|data~93_combout ;
wire	\macro_inst|controller|sm_pwm|data~94_combout ;
wire	\macro_inst|controller|sm_pwm|data~95_combout ;
wire	\macro_inst|controller|sm_pwm|data~96_combout ;
wire	\macro_inst|controller|sm_pwm|data~97_combout ;
wire	\macro_inst|controller|sm_pwm|data~98_combout ;
wire	\macro_inst|controller|sm_pwm|data~99_combout ;
wire	\macro_inst|controller|sm_pwm|data~9_combout ;
wire	[15:0] \macro_inst|controller|sm_pwm|motor_flags ;
//wire	\macro_inst|controller|sm_pwm|motor_flags [0];
wire	\macro_inst|controller|sm_pwm|motor_flags[0]~0_combout ;
wire	\macro_inst|controller|sm_pwm|motor_flags[0]~1_combout ;
wire	\macro_inst|controller|sm_pwm|motor_flags[0]~2_combout ;
wire	\macro_inst|controller|sm_pwm|motor_flags[0]~3_combout ;
wire	\macro_inst|controller|sm_pwm|motor_flags[0]~4_combout ;
wire	\macro_inst|controller|sm_pwm|motor_flags[0]~5_combout ;
wire	\macro_inst|controller|sm_pwm|motor_flags[0]~6_combout ;
wire	\macro_inst|controller|sm_pwm|motor_flags[0]~7_combout ;
//wire	\macro_inst|controller|sm_pwm|motor_flags [10];
//wire	\macro_inst|controller|sm_pwm|motor_flags [11];
//wire	\macro_inst|controller|sm_pwm|motor_flags [12];
//wire	\macro_inst|controller|sm_pwm|motor_flags [13];
//wire	\macro_inst|controller|sm_pwm|motor_flags [14];
//wire	\macro_inst|controller|sm_pwm|motor_flags [15];
//wire	\macro_inst|controller|sm_pwm|motor_flags [1];
//wire	\macro_inst|controller|sm_pwm|motor_flags [2];
//wire	\macro_inst|controller|sm_pwm|motor_flags [3];
//wire	\macro_inst|controller|sm_pwm|motor_flags [4];
//wire	\macro_inst|controller|sm_pwm|motor_flags [5];
//wire	\macro_inst|controller|sm_pwm|motor_flags [6];
//wire	\macro_inst|controller|sm_pwm|motor_flags [7];
//wire	\macro_inst|controller|sm_pwm|motor_flags [8];
//wire	\macro_inst|controller|sm_pwm|motor_flags [9];
wire	[7:0] \macro_inst|controller|sm_pwm|pwmCnt ;
//wire	\macro_inst|controller|sm_pwm|pwmCnt [0];
//wire	\macro_inst|controller|sm_pwm|pwmCnt [1];
//wire	\macro_inst|controller|sm_pwm|pwmCnt [2];
//wire	\macro_inst|controller|sm_pwm|pwmCnt [3];
//wire	\macro_inst|controller|sm_pwm|pwmCnt [4];
//wire	\macro_inst|controller|sm_pwm|pwmCnt [5];
//wire	\macro_inst|controller|sm_pwm|pwmCnt [6];
//wire	\macro_inst|controller|sm_pwm|pwmCnt [7];
wire	\macro_inst|controller|sm_pwm|pwmCnt~0_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][0]~49_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][5]~48_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[0][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][0]~87_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][5]~86_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][8]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[10][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][0]~39_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][5]~38_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[11][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][0]~89_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][5]~88_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[12][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][0]~41_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][5]~40_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[13][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][0]~91_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][5]~90_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[14][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][0]~43_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][5]~42_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[15][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][0]~93_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][5]~92_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[16][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][0]~45_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][15]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][5]~44_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[17][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][0]~95_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][5]~94_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[18][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][0]~47_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][15]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][5]~46_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[19][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][0]~1_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][5]~0_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[1][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][0]~53_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][15]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][5]~52_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[20][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][0]~5_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][5]~4_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[21][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][0]~55_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][5]~54_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[22][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][0]~7_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][5]~6_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[23][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][0]~57_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][5]~56_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[24][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][0]~9_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][5]~8_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[25][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][0]~59_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][5]~58_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[26][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][0]~11_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][10]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][11]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][12]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][13]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][5]~10_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[27][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][0]~61_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][5]~60_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[28][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][0]~13_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][5]~12_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[29][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][0]~51_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][12]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][5]~50_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[2][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][0]~63_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][5]~62_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[30][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][0]~15_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][5]~14_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[31][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][0]~65_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][5]~64_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[32][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][0]~17_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][5]~16_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][8]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[33][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][0]~67_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][12]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][1]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][3]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][5]~66_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[34][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][0]~19_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][15]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][5]~18_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[35][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][0]~69_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][5]~68_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[36][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][0]~21_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][5]~20_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[37][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][0]~71_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][5]~70_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[38][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][0]~23_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][5]~22_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[39][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][0]~3_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][10]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][13]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][5]~2_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[3][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][0]~75_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][5]~74_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[40][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][0]~27_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][5]~26_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[41][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][0]~77_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][5]~76_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[42][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][0]~29_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][15]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][5]~28_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[43][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][0]~79_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][5]~78_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[44][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][0]~31_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][15]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][5]~30_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[45][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][0]~81_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][15]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][5]~80_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[46][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][0]~33_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][5]~32_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[47][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][0]~73_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][5]~72_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[4][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][0]~25_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][15]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][5]~24_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[5][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][0]~83_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][5]~82_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[6][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][0]~35_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][15]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][5]~34_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[7][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][0]~85_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][5]~84_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[8][9]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][0]~37_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][0]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][10]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][11]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][12]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][13]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][14]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][15]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][15]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][1]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][2]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][3]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][4]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][5]~36_combout ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][5]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][6]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][7]__feeder__LutOut ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][7]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][8]~q ;
wire	\macro_inst|controller|sm_pwm|pwmList[9][9]~q ;
wire	\macro_inst|mem_ahb_hrdata[0]~0_combout ;
wire	\macro_inst|mem_ahb_hrdata[10]~10_combout ;
wire	\macro_inst|mem_ahb_hrdata[11]~11_combout ;
wire	\macro_inst|mem_ahb_hrdata[12]~12_combout ;
wire	\macro_inst|mem_ahb_hrdata[13]~13_combout ;
wire	\macro_inst|mem_ahb_hrdata[14]~14_combout ;
wire	\macro_inst|mem_ahb_hrdata[15]~15_combout ;
wire	\macro_inst|mem_ahb_hrdata[16]~16_combout ;
wire	\macro_inst|mem_ahb_hrdata[17]~17_combout ;
wire	\macro_inst|mem_ahb_hrdata[18]~18_combout ;
wire	\macro_inst|mem_ahb_hrdata[19]~19_combout ;
wire	\macro_inst|mem_ahb_hrdata[1]~1_combout ;
wire	\macro_inst|mem_ahb_hrdata[20]~20_combout ;
wire	\macro_inst|mem_ahb_hrdata[21]~21_combout ;
wire	\macro_inst|mem_ahb_hrdata[22]~22_combout ;
wire	\macro_inst|mem_ahb_hrdata[23]~23_combout ;
wire	\macro_inst|mem_ahb_hrdata[24]~24_combout ;
wire	\macro_inst|mem_ahb_hrdata[25]~25_combout ;
wire	\macro_inst|mem_ahb_hrdata[26]~26_combout ;
wire	\macro_inst|mem_ahb_hrdata[27]~27_combout ;
wire	\macro_inst|mem_ahb_hrdata[28]~28_combout ;
wire	\macro_inst|mem_ahb_hrdata[29]~29_combout ;
wire	\macro_inst|mem_ahb_hrdata[2]~2_combout ;
wire	\macro_inst|mem_ahb_hrdata[30]~30_combout ;
wire	\macro_inst|mem_ahb_hrdata[31]~31_combout ;
wire	\macro_inst|mem_ahb_hrdata[3]~3_combout ;
wire	\macro_inst|mem_ahb_hrdata[4]~4_combout ;
wire	\macro_inst|mem_ahb_hrdata[5]~5_combout ;
wire	\macro_inst|mem_ahb_hrdata[6]~6_combout ;
wire	\macro_inst|mem_ahb_hrdata[7]~7_combout ;
wire	\macro_inst|mem_ahb_hrdata[8]~8_combout ;
wire	\macro_inst|mem_ahb_hrdata[9]~9_combout ;
wire	\macro_inst|serial_lim_input_inst|Add1~0_combout ;
wire	\macro_inst|serial_lim_input_inst|Decoder0~0_combout ;
wire	\macro_inst|serial_lim_input_inst|Decoder0~1_combout ;
wire	\macro_inst|serial_lim_input_inst|Decoder0~2_combout ;
wire	\macro_inst|serial_lim_input_inst|Decoder0~3_combout ;
wire	\macro_inst|serial_lim_input_inst|Decoder0~4_combout ;
wire	\macro_inst|serial_lim_input_inst|Decoder0~5_combout ;
wire	\macro_inst|serial_lim_input_inst|Decoder0~6_combout ;
wire	\macro_inst|serial_lim_input_inst|Decoder0~7_combout ;
wire	\macro_inst|serial_lim_input_inst|Decoder0~8_combout ;
wire	\macro_inst|serial_lim_input_inst|Equal0~0_combout ;
wire	\macro_inst|serial_lim_input_inst|Equal0~1_combout ;
wire	\macro_inst|serial_lim_input_inst|Equal0~2_combout ;
wire	\macro_inst|serial_lim_input_inst|Equal0~3_combout ;
wire	\macro_inst|serial_lim_input_inst|Equal0~4_combout ;
wire	\macro_inst|serial_lim_input_inst|Equal2~0_combout ;
wire	\macro_inst|serial_lim_input_inst|Equal2~1_combout ;
wire	\macro_inst|serial_lim_input_inst|Equal2~2_combout ;
wire	\macro_inst|serial_lim_input_inst|Equal2~3_combout ;
wire	\macro_inst|serial_lim_input_inst|Equal2~4_combout ;
wire	\macro_inst|serial_lim_input_inst|Selector18~0_combout ;
wire	\macro_inst|serial_lim_input_inst|Selector19~0_combout ;
wire	\macro_inst|serial_lim_input_inst|Selector20~2_combout ;
wire	\macro_inst|serial_lim_input_inst|Selector20~3_combout ;
wire	\macro_inst|serial_lim_input_inst|Selector20~4_combout ;
wire	\macro_inst|serial_lim_input_inst|Selector20~5_combout ;
wire	\macro_inst|serial_lim_input_inst|ahb_read_transfer~combout ;
wire	[2:0] \macro_inst|serial_lim_input_inst|bit_counter ;
//wire	\macro_inst|serial_lim_input_inst|bit_counter [0];
wire	\macro_inst|serial_lim_input_inst|bit_counter[0]~4_combout ;
//wire	\macro_inst|serial_lim_input_inst|bit_counter [1];
wire	\macro_inst|serial_lim_input_inst|bit_counter[1]~0_combout ;
wire	\macro_inst|serial_lim_input_inst|bit_counter[1]~1_combout ;
wire	\macro_inst|serial_lim_input_inst|bit_counter[1]~3_combout ;
//wire	\macro_inst|serial_lim_input_inst|bit_counter [2];
wire	\macro_inst|serial_lim_input_inst|bit_counter[2]~2_combout ;
wire	\macro_inst|serial_lim_input_inst|capture_done~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|capture_done~q ;
wire	[47:0] \macro_inst|serial_lim_input_inst|captured_data ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [0];
wire	\macro_inst|serial_lim_input_inst|captured_data[0]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [10];
wire	\macro_inst|serial_lim_input_inst|captured_data[10]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [11];
wire	\macro_inst|serial_lim_input_inst|captured_data[11]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [12];
wire	\macro_inst|serial_lim_input_inst|captured_data[12]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [13];
wire	\macro_inst|serial_lim_input_inst|captured_data[13]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [14];
wire	\macro_inst|serial_lim_input_inst|captured_data[14]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [15];
wire	\macro_inst|serial_lim_input_inst|captured_data[15]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [16];
//wire	\macro_inst|serial_lim_input_inst|captured_data [17];
wire	\macro_inst|serial_lim_input_inst|captured_data[17]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [18];
wire	\macro_inst|serial_lim_input_inst|captured_data[18]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [19];
wire	\macro_inst|serial_lim_input_inst|captured_data[19]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [1];
wire	\macro_inst|serial_lim_input_inst|captured_data[1]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [20];
wire	\macro_inst|serial_lim_input_inst|captured_data[20]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [21];
wire	\macro_inst|serial_lim_input_inst|captured_data[21]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [22];
wire	\macro_inst|serial_lim_input_inst|captured_data[22]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [23];
wire	\macro_inst|serial_lim_input_inst|captured_data[23]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [24];
wire	\macro_inst|serial_lim_input_inst|captured_data[24]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [25];
wire	\macro_inst|serial_lim_input_inst|captured_data[25]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [26];
wire	\macro_inst|serial_lim_input_inst|captured_data[26]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [27];
wire	\macro_inst|serial_lim_input_inst|captured_data[27]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [28];
wire	\macro_inst|serial_lim_input_inst|captured_data[28]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [29];
wire	\macro_inst|serial_lim_input_inst|captured_data[29]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [2];
wire	\macro_inst|serial_lim_input_inst|captured_data[2]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [30];
wire	\macro_inst|serial_lim_input_inst|captured_data[30]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [31];
wire	\macro_inst|serial_lim_input_inst|captured_data[31]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [32];
wire	\macro_inst|serial_lim_input_inst|captured_data[32]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [33];
wire	\macro_inst|serial_lim_input_inst|captured_data[33]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [34];
wire	\macro_inst|serial_lim_input_inst|captured_data[34]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [35];
wire	\macro_inst|serial_lim_input_inst|captured_data[35]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [36];
//wire	\macro_inst|serial_lim_input_inst|captured_data [37];
wire	\macro_inst|serial_lim_input_inst|captured_data[37]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [38];
wire	\macro_inst|serial_lim_input_inst|captured_data[38]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [39];
wire	\macro_inst|serial_lim_input_inst|captured_data[39]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [3];
wire	\macro_inst|serial_lim_input_inst|captured_data[3]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [40];
wire	\macro_inst|serial_lim_input_inst|captured_data[40]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [41];
wire	\macro_inst|serial_lim_input_inst|captured_data[41]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [42];
wire	\macro_inst|serial_lim_input_inst|captured_data[42]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [43];
wire	\macro_inst|serial_lim_input_inst|captured_data[43]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [44];
wire	\macro_inst|serial_lim_input_inst|captured_data[44]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [45];
wire	\macro_inst|serial_lim_input_inst|captured_data[45]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [46];
wire	\macro_inst|serial_lim_input_inst|captured_data[46]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [47];
wire	\macro_inst|serial_lim_input_inst|captured_data[47]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [4];
//wire	\macro_inst|serial_lim_input_inst|captured_data [5];
wire	\macro_inst|serial_lim_input_inst|captured_data[5]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [6];
wire	\macro_inst|serial_lim_input_inst|captured_data[6]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [7];
wire	\macro_inst|serial_lim_input_inst|captured_data[7]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [8];
wire	\macro_inst|serial_lim_input_inst|captured_data[8]~feeder_combout ;
//wire	\macro_inst|serial_lim_input_inst|captured_data [9];
wire	[15:0] \macro_inst|serial_lim_input_inst|load_counter ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [0];
wire	\macro_inst|serial_lim_input_inst|load_counter[0]~17_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[0]~18 ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [10];
wire	\macro_inst|serial_lim_input_inst|load_counter[10]~38_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[10]~39 ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [11];
wire	\macro_inst|serial_lim_input_inst|load_counter[11]~40_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[11]~41 ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [12];
wire	\macro_inst|serial_lim_input_inst|load_counter[12]~42_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[12]~43 ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [13];
wire	\macro_inst|serial_lim_input_inst|load_counter[13]~44_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[13]~45 ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [14];
wire	\macro_inst|serial_lim_input_inst|load_counter[14]~16_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[14]~19_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[14]~46_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[14]~47 ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [15];
wire	\macro_inst|serial_lim_input_inst|load_counter[15]~48_combout ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [1];
wire	\macro_inst|serial_lim_input_inst|load_counter[1]~20_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[1]~21 ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [2];
wire	\macro_inst|serial_lim_input_inst|load_counter[2]~22_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[2]~23 ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [3];
wire	\macro_inst|serial_lim_input_inst|load_counter[3]~24_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[3]~25 ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [4];
wire	\macro_inst|serial_lim_input_inst|load_counter[4]~26_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[4]~27 ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [5];
wire	\macro_inst|serial_lim_input_inst|load_counter[5]~28_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[5]~29 ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [6];
wire	\macro_inst|serial_lim_input_inst|load_counter[6]~30_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[6]~31 ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [7];
wire	\macro_inst|serial_lim_input_inst|load_counter[7]~32_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[7]~33 ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [8];
wire	\macro_inst|serial_lim_input_inst|load_counter[8]~34_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[8]~35 ;
//wire	\macro_inst|serial_lim_input_inst|load_counter [9];
wire	\macro_inst|serial_lim_input_inst|load_counter[9]~36_combout ;
wire	\macro_inst|serial_lim_input_inst|load_counter[9]~37 ;
wire	\macro_inst|serial_lim_input_inst|load~0_combout ;
wire	\macro_inst|serial_lim_input_inst|load~1_combout ;
wire	\macro_inst|serial_lim_input_inst|load~q ;
wire	[31:0] \macro_inst|serial_lim_input_inst|mem_ahb_hrdata ;
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [0];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [10];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [11];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [12];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [13];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [14];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [15];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [16];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [17];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [18];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [19];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [1];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [20];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [21];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [22];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [23];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [24];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [25];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [26];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [27];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [28];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [29];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [2];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [30];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [31];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [3];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [4];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [5];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [6];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [7];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [8];
//wire	\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [9];
wire	\macro_inst|serial_lim_input_inst|read_chunk[0]~0_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[10]~10_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[11]~11_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[12]~12_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[13]~13_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[14]~14_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[15]~15_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[16]~16_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[17]~17_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[18]~18_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[19]~19_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[1]~1_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[20]~20_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[21]~21_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[22]~22_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[23]~23_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[24]~24_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[25]~25_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[26]~26_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[27]~27_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[28]~28_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[29]~29_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[2]~2_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[30]~30_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[31]~31_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[3]~3_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[4]~4_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[5]~5_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[6]~6_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[7]~7_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[8]~8_combout ;
wire	\macro_inst|serial_lim_input_inst|read_chunk[9]~9_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][0]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][0]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][1]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][1]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][2]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][2]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][3]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][3]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][4]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][5]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][5]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][6]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][6]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][7]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[0][7]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][0]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][0]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][1]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][1]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][2]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][2]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][3]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][3]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][4]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][4]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][5]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][5]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][6]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][6]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][7]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[1][7]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[2][0]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[2][1]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[2][1]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[2][2]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[2][3]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[2][3]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[2][4]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[2][4]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[2][5]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[2][5]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[2][6]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[2][7]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[2][7]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[3][0]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[3][0]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[3][1]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[3][2]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[3][2]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[3][3]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[3][4]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[3][4]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[3][5]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[3][6]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[3][6]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[3][7]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][0]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][1]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][1]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][2]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][2]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][3]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][3]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][4]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][4]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][5]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][5]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][6]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][6]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][7]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[4][7]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[5][0]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[5][0]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[5][1]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[5][1]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[5][2]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[5][3]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[5][3]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[5][4]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[5][4]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[5][5]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[5][5]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[5][6]~q ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[5][7]~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_buffer[5][7]~q ;
wire	[15:0] \macro_inst|serial_lim_input_inst|shift_div_counter ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [0];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[0]~16_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[0]~17 ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [10];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[10]~37_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[10]~38 ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [11];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[11]~39_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[11]~40 ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [12];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[12]~41_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[12]~42 ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [13];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[13]~43_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[13]~44 ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [14];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[14]~45_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[14]~46 ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [15];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[15]~47_combout ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [1];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[1]~18_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[1]~19 ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [2];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[2]~21_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[2]~22 ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [3];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[3]~23_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[3]~24 ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [4];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[4]~25_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[4]~26 ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [5];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[5]~27_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[5]~28 ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [6];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[6]~29_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[6]~30 ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [7];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[7]~31_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[7]~32 ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [8];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[8]~33_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[8]~34 ;
//wire	\macro_inst|serial_lim_input_inst|shift_div_counter [9];
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[9]~35_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_div_counter[9]~36 ;
wire	\macro_inst|serial_lim_input_inst|shift_enable~0_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_enable~1_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_enable~2_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_enable~q ;
wire	\macro_inst|serial_lim_input_inst|shift_out_d~q ;
wire	\macro_inst|serial_lim_input_inst|shift_out~0_combout ;
wire	\macro_inst|serial_lim_input_inst|shift_out~q ;
wire	\macro_inst|serial_lim_input_inst|shift_rise~combout ;
wire	\macro_inst|serial_lim_input_inst|shift~combout ;
wire	\macro_inst|serial_lim_input_inst|state_reg.STATE_IDLE~q ;
wire	\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q ;
wire	\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ;
wire	\macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT~q ;
wire	\macro_inst|serial_lim_input_inst|trigger_sync0~q ;
wire	\macro_inst|serial_lim_input_inst|trigger_sync1~feeder_combout ;
wire	\macro_inst|serial_lim_input_inst|trigger_sync1~q ;
wire	[4:0] \pll_inst|auto_generated|clk ;
//wire	\pll_inst|auto_generated|clk [0];
//wire	\pll_inst|auto_generated|clk [1];
//wire	\pll_inst|auto_generated|clk [2];
//wire	\pll_inst|auto_generated|clk [3];
//wire	\pll_inst|auto_generated|clk [4];
wire	[4:0] \pll_inst|auto_generated|pll1_CLK_bus ;
//wire	\pll_inst|auto_generated|pll1_CLK_bus [0];
//wire	\pll_inst|auto_generated|pll1_CLK_bus [1];
//wire	\pll_inst|auto_generated|pll1_CLK_bus [2];
//wire	\pll_inst|auto_generated|pll1_CLK_bus [3];
//wire	\pll_inst|auto_generated|pll1_CLK_bus [4];
wire	\pll_inst|auto_generated|pll1~FBOUT ;
wire	\pll_inst|auto_generated|pll_lock_sync~feeder_combout ;
wire	\pll_inst|auto_generated|pll_lock_sync~q ;
wire	\rv32.dmactive ;
wire	\rv32.ext_dma_DMACCLR[0] ;
wire	\rv32.ext_dma_DMACCLR[1] ;
wire	\rv32.ext_dma_DMACCLR[2] ;
wire	\rv32.ext_dma_DMACCLR[3] ;
wire	\rv32.ext_dma_DMACTC[0] ;
wire	\rv32.ext_dma_DMACTC[1] ;
wire	\rv32.ext_dma_DMACTC[2] ;
wire	\rv32.ext_dma_DMACTC[3] ;
wire	\rv32.gpio0_io_out_data[0] ;
wire	\rv32.gpio0_io_out_data[1] ;
wire	\rv32.gpio0_io_out_data[2] ;
wire	\rv32.gpio0_io_out_data[3] ;
wire	\rv32.gpio0_io_out_data[4] ;
wire	\rv32.gpio0_io_out_data[5] ;
wire	\rv32.gpio0_io_out_data[6] ;
wire	\rv32.gpio0_io_out_data[7] ;
wire	\rv32.gpio0_io_out_en[0] ;
wire	\rv32.gpio0_io_out_en[1] ;
wire	\rv32.gpio0_io_out_en[2] ;
wire	\rv32.gpio0_io_out_en[3] ;
wire	\rv32.gpio0_io_out_en[4] ;
wire	\rv32.gpio0_io_out_en[5] ;
wire	\rv32.gpio0_io_out_en[6] ;
wire	\rv32.gpio0_io_out_en[7] ;
wire	\rv32.gpio1_io_out_data[0] ;
wire	\rv32.gpio1_io_out_data[1] ;
wire	\rv32.gpio1_io_out_data[2] ;
wire	\rv32.gpio1_io_out_data[3] ;
wire	\rv32.gpio1_io_out_data[4] ;
wire	\rv32.gpio1_io_out_data[5] ;
wire	\rv32.gpio1_io_out_data[6] ;
wire	\rv32.gpio1_io_out_data[7] ;
wire	\rv32.gpio1_io_out_en[0] ;
wire	\rv32.gpio1_io_out_en[1] ;
wire	\rv32.gpio1_io_out_en[2] ;
wire	\rv32.gpio1_io_out_en[3] ;
wire	\rv32.gpio1_io_out_en[4] ;
wire	\rv32.gpio1_io_out_en[5] ;
wire	\rv32.gpio1_io_out_en[6] ;
wire	\rv32.gpio1_io_out_en[7] ;
wire	\rv32.gpio2_io_out_data[0] ;
wire	\rv32.gpio2_io_out_data[1] ;
wire	\rv32.gpio2_io_out_data[2] ;
wire	\rv32.gpio2_io_out_data[3] ;
wire	\rv32.gpio2_io_out_data[4] ;
wire	\rv32.gpio2_io_out_data[5] ;
wire	\rv32.gpio2_io_out_data[6] ;
wire	\rv32.gpio2_io_out_data[7] ;
wire	\rv32.gpio2_io_out_en[0] ;
wire	\rv32.gpio2_io_out_en[1] ;
wire	\rv32.gpio2_io_out_en[2] ;
wire	\rv32.gpio2_io_out_en[3] ;
wire	\rv32.gpio2_io_out_en[4] ;
wire	\rv32.gpio2_io_out_en[5] ;
wire	\rv32.gpio2_io_out_en[6] ;
wire	\rv32.gpio2_io_out_en[7] ;
wire	\rv32.gpio3_io_out_data[0] ;
wire	\rv32.gpio3_io_out_data[1] ;
wire	\rv32.gpio3_io_out_data[2] ;
wire	\rv32.gpio3_io_out_data[3] ;
wire	\rv32.gpio3_io_out_data[4] ;
wire	\rv32.gpio3_io_out_data[5] ;
wire	\rv32.gpio3_io_out_data[6] ;
wire	\rv32.gpio3_io_out_data[7] ;
wire	\rv32.gpio3_io_out_en[0] ;
wire	\rv32.gpio3_io_out_en[1] ;
wire	\rv32.gpio3_io_out_en[2] ;
wire	\rv32.gpio3_io_out_en[3] ;
wire	\rv32.gpio3_io_out_en[4] ;
wire	\rv32.gpio3_io_out_en[5] ;
wire	\rv32.gpio3_io_out_en[6] ;
wire	\rv32.gpio3_io_out_en[7] ;
wire	\rv32.gpio4_io_out_data[0] ;
wire	\rv32.gpio4_io_out_data[1] ;
wire	\rv32.gpio4_io_out_data[2] ;
wire	\rv32.gpio4_io_out_data[3] ;
wire	\rv32.gpio4_io_out_data[4] ;
wire	\rv32.gpio4_io_out_data[5] ;
wire	\rv32.gpio4_io_out_data[6] ;
wire	\rv32.gpio4_io_out_data[7] ;
wire	\rv32.gpio4_io_out_en[0] ;
wire	\rv32.gpio4_io_out_en[1] ;
wire	\rv32.gpio4_io_out_en[2] ;
wire	\rv32.gpio4_io_out_en[3] ;
wire	\rv32.gpio4_io_out_en[4] ;
wire	\rv32.gpio4_io_out_en[5] ;
wire	\rv32.gpio4_io_out_en[6] ;
wire	\rv32.gpio4_io_out_en[7] ;
wire	\rv32.gpio5_io_out_data[0] ;
wire	\rv32.gpio5_io_out_data[1] ;
wire	\rv32.gpio5_io_out_data[2] ;
wire	\rv32.gpio5_io_out_data[3] ;
wire	\rv32.gpio5_io_out_data[4] ;
wire	\rv32.gpio5_io_out_data[5] ;
wire	\rv32.gpio5_io_out_data[6] ;
wire	\rv32.gpio5_io_out_data[7] ;
wire	\rv32.gpio5_io_out_en[0] ;
wire	\rv32.gpio5_io_out_en[1] ;
wire	\rv32.gpio5_io_out_en[2] ;
wire	\rv32.gpio5_io_out_en[3] ;
wire	\rv32.gpio5_io_out_en[4] ;
wire	\rv32.gpio5_io_out_en[5] ;
wire	\rv32.gpio5_io_out_en[6] ;
wire	\rv32.gpio5_io_out_en[7] ;
wire	\rv32.gpio6_io_out_data[0] ;
wire	\rv32.gpio6_io_out_data[1] ;
wire	\rv32.gpio6_io_out_data[2] ;
wire	\rv32.gpio6_io_out_data[3] ;
wire	\rv32.gpio6_io_out_data[4] ;
wire	\rv32.gpio6_io_out_data[5] ;
wire	\rv32.gpio6_io_out_data[6] ;
wire	\rv32.gpio6_io_out_data[7] ;
wire	\rv32.gpio6_io_out_en[0] ;
wire	\rv32.gpio6_io_out_en[1] ;
wire	\rv32.gpio6_io_out_en[2] ;
wire	\rv32.gpio6_io_out_en[3] ;
wire	\rv32.gpio6_io_out_en[4] ;
wire	\rv32.gpio6_io_out_en[5] ;
wire	\rv32.gpio6_io_out_en[6] ;
wire	\rv32.gpio6_io_out_en[7] ;
wire	\rv32.gpio7_io_out_data[0] ;
wire	\rv32.gpio7_io_out_data[1] ;
wire	\rv32.gpio7_io_out_data[2] ;
wire	\rv32.gpio7_io_out_data[3] ;
wire	\rv32.gpio7_io_out_data[4] ;
wire	\rv32.gpio7_io_out_data[5] ;
wire	\rv32.gpio7_io_out_data[6] ;
wire	\rv32.gpio7_io_out_data[7] ;
wire	\rv32.gpio7_io_out_en[0] ;
wire	\rv32.gpio7_io_out_en[1] ;
wire	\rv32.gpio7_io_out_en[2] ;
wire	\rv32.gpio7_io_out_en[3] ;
wire	\rv32.gpio7_io_out_en[4] ;
wire	\rv32.gpio7_io_out_en[5] ;
wire	\rv32.gpio7_io_out_en[6] ;
wire	\rv32.gpio7_io_out_en[7] ;
wire	\rv32.gpio8_io_out_data[0] ;
wire	\rv32.gpio8_io_out_data[1] ;
wire	\rv32.gpio8_io_out_data[2] ;
wire	\rv32.gpio8_io_out_data[3] ;
wire	\rv32.gpio8_io_out_data[4] ;
wire	\rv32.gpio8_io_out_data[5] ;
wire	\rv32.gpio8_io_out_data[6] ;
wire	\rv32.gpio8_io_out_data[7] ;
wire	\rv32.gpio8_io_out_en[0] ;
wire	\rv32.gpio8_io_out_en[1] ;
wire	\rv32.gpio8_io_out_en[2] ;
wire	\rv32.gpio8_io_out_en[3] ;
wire	\rv32.gpio8_io_out_en[4] ;
wire	\rv32.gpio8_io_out_en[5] ;
wire	\rv32.gpio8_io_out_en[6] ;
wire	\rv32.gpio8_io_out_en[7] ;
wire	\rv32.gpio9_io_out_data[0] ;
wire	\rv32.gpio9_io_out_data[1] ;
wire	\rv32.gpio9_io_out_data[2] ;
wire	\rv32.gpio9_io_out_data[3] ;
wire	\rv32.gpio9_io_out_data[4] ;
wire	\rv32.gpio9_io_out_data[5] ;
wire	\rv32.gpio9_io_out_data[6] ;
wire	\rv32.gpio9_io_out_data[7] ;
wire	\rv32.gpio9_io_out_en[0] ;
wire	\rv32.gpio9_io_out_en[1] ;
wire	\rv32.gpio9_io_out_en[2] ;
wire	\rv32.gpio9_io_out_en[3] ;
wire	\rv32.gpio9_io_out_en[4] ;
wire	\rv32.gpio9_io_out_en[5] ;
wire	\rv32.gpio9_io_out_en[6] ;
wire	\rv32.gpio9_io_out_en[7] ;
wire	\rv32.mem_ahb_haddr[0] ;
wire	\rv32.mem_ahb_haddr[10] ;
wire	\rv32.mem_ahb_haddr[11] ;
wire	\rv32.mem_ahb_haddr[12] ;
wire	\rv32.mem_ahb_haddr[13] ;
wire	\rv32.mem_ahb_haddr[14] ;
wire	\rv32.mem_ahb_haddr[15] ;
wire	\rv32.mem_ahb_haddr[16] ;
wire	\rv32.mem_ahb_haddr[17] ;
wire	\rv32.mem_ahb_haddr[18] ;
wire	\rv32.mem_ahb_haddr[19] ;
wire	\rv32.mem_ahb_haddr[1] ;
wire	\rv32.mem_ahb_haddr[20] ;
wire	\rv32.mem_ahb_haddr[21] ;
wire	\rv32.mem_ahb_haddr[22] ;
wire	\rv32.mem_ahb_haddr[23] ;
wire	\rv32.mem_ahb_haddr[24] ;
wire	\rv32.mem_ahb_haddr[25] ;
wire	\rv32.mem_ahb_haddr[26] ;
wire	\rv32.mem_ahb_haddr[27] ;
wire	\rv32.mem_ahb_haddr[28] ;
wire	\rv32.mem_ahb_haddr[29] ;
wire	\rv32.mem_ahb_haddr[2] ;
wire	\rv32.mem_ahb_haddr[30] ;
wire	\rv32.mem_ahb_haddr[31] ;
wire	\rv32.mem_ahb_haddr[3] ;
wire	\rv32.mem_ahb_haddr[3]__SyncReset_X56_Y3_SIG ;
wire	\rv32.mem_ahb_haddr[3]__SyncReset_X56_Y5_SIG ;
wire	\rv32.mem_ahb_haddr[3]__SyncReset_X57_Y5_SIG ;
wire	\rv32.mem_ahb_haddr[4] ;
wire	\rv32.mem_ahb_haddr[5] ;
wire	\rv32.mem_ahb_haddr[6] ;
wire	\rv32.mem_ahb_haddr[7] ;
wire	\rv32.mem_ahb_haddr[8] ;
wire	\rv32.mem_ahb_haddr[9] ;
wire	\rv32.mem_ahb_hburst[0] ;
wire	\rv32.mem_ahb_hburst[1] ;
wire	\rv32.mem_ahb_hburst[2] ;
wire	\rv32.mem_ahb_hready ;
wire	\rv32.mem_ahb_hsize[0] ;
wire	\rv32.mem_ahb_hsize[1] ;
wire	\rv32.mem_ahb_hsize[2] ;
wire	\rv32.mem_ahb_htrans[0] ;
wire	\rv32.mem_ahb_htrans[1] ;
wire	\rv32.mem_ahb_hwdata[0] ;
wire	\rv32.mem_ahb_hwdata[10] ;
wire	\rv32.mem_ahb_hwdata[11] ;
wire	\rv32.mem_ahb_hwdata[12] ;
wire	\rv32.mem_ahb_hwdata[13] ;
wire	\rv32.mem_ahb_hwdata[14] ;
wire	\rv32.mem_ahb_hwdata[15] ;
wire	\rv32.mem_ahb_hwdata[16] ;
wire	\rv32.mem_ahb_hwdata[17] ;
wire	\rv32.mem_ahb_hwdata[18] ;
wire	\rv32.mem_ahb_hwdata[19] ;
wire	\rv32.mem_ahb_hwdata[1] ;
wire	\rv32.mem_ahb_hwdata[20] ;
wire	\rv32.mem_ahb_hwdata[21] ;
wire	\rv32.mem_ahb_hwdata[22] ;
wire	\rv32.mem_ahb_hwdata[23] ;
wire	\rv32.mem_ahb_hwdata[24] ;
wire	\rv32.mem_ahb_hwdata[25] ;
wire	\rv32.mem_ahb_hwdata[26] ;
wire	\rv32.mem_ahb_hwdata[27] ;
wire	\rv32.mem_ahb_hwdata[28] ;
wire	\rv32.mem_ahb_hwdata[29] ;
wire	\rv32.mem_ahb_hwdata[2] ;
wire	\rv32.mem_ahb_hwdata[30] ;
wire	\rv32.mem_ahb_hwdata[31] ;
wire	\rv32.mem_ahb_hwdata[3] ;
wire	\rv32.mem_ahb_hwdata[4] ;
wire	\rv32.mem_ahb_hwdata[5] ;
wire	\rv32.mem_ahb_hwdata[6] ;
wire	\rv32.mem_ahb_hwdata[7] ;
wire	\rv32.mem_ahb_hwdata[8] ;
wire	\rv32.mem_ahb_hwdata[9] ;
wire	\rv32.mem_ahb_hwrite ;
wire	\rv32.resetn_out ;
wire	\rv32.slave_ahb_hrdata[0] ;
wire	\rv32.slave_ahb_hrdata[10] ;
wire	\rv32.slave_ahb_hrdata[11] ;
wire	\rv32.slave_ahb_hrdata[12] ;
wire	\rv32.slave_ahb_hrdata[13] ;
wire	\rv32.slave_ahb_hrdata[14] ;
wire	\rv32.slave_ahb_hrdata[15] ;
wire	\rv32.slave_ahb_hrdata[16] ;
wire	\rv32.slave_ahb_hrdata[17] ;
wire	\rv32.slave_ahb_hrdata[18] ;
wire	\rv32.slave_ahb_hrdata[19] ;
wire	\rv32.slave_ahb_hrdata[1] ;
wire	\rv32.slave_ahb_hrdata[20] ;
wire	\rv32.slave_ahb_hrdata[21] ;
wire	\rv32.slave_ahb_hrdata[22] ;
wire	\rv32.slave_ahb_hrdata[23] ;
wire	\rv32.slave_ahb_hrdata[24] ;
wire	\rv32.slave_ahb_hrdata[25] ;
wire	\rv32.slave_ahb_hrdata[26] ;
wire	\rv32.slave_ahb_hrdata[27] ;
wire	\rv32.slave_ahb_hrdata[28] ;
wire	\rv32.slave_ahb_hrdata[29] ;
wire	\rv32.slave_ahb_hrdata[2] ;
wire	\rv32.slave_ahb_hrdata[30] ;
wire	\rv32.slave_ahb_hrdata[31] ;
wire	\rv32.slave_ahb_hrdata[3] ;
wire	\rv32.slave_ahb_hrdata[4] ;
wire	\rv32.slave_ahb_hrdata[5] ;
wire	\rv32.slave_ahb_hrdata[6] ;
wire	\rv32.slave_ahb_hrdata[7] ;
wire	\rv32.slave_ahb_hrdata[8] ;
wire	\rv32.slave_ahb_hrdata[9] ;
wire	\rv32.slave_ahb_hreadyout ;
wire	\rv32.slave_ahb_hresp ;
wire	\rv32.swj_JTAGIR[0] ;
wire	\rv32.swj_JTAGIR[1] ;
wire	\rv32.swj_JTAGIR[2] ;
wire	\rv32.swj_JTAGIR[3] ;
wire	\rv32.swj_JTAGNSW ;
wire	\rv32.swj_JTAGSTATE[0] ;
wire	\rv32.swj_JTAGSTATE[1] ;
wire	\rv32.swj_JTAGSTATE[2] ;
wire	\rv32.swj_JTAGSTATE[3] ;
wire	\rv32.sys_ctrl_clkSource[0] ;
wire	\rv32.sys_ctrl_clkSource[1] ;
wire	\rv32.sys_ctrl_hseBypass ;
wire	\rv32.sys_ctrl_hseEnable ;
wire	\rv32.sys_ctrl_pllEnable ;
wire	\rv32.sys_ctrl_sleep ;
wire	\rv32.sys_ctrl_standby ;
wire	\rv32.sys_ctrl_stop ;
wire	\sys_resetn~clkctrl_outclk ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y3_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X47_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X47_Y3_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y3_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y1_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y4_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y1_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y4_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y1_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y3_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y9_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y12_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y1_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y3_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y5_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y6_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y8_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y10_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y12_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y3_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y4_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y5_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y7_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y8_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y11_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y3_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y4_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y6_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y3_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y7_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y10_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y1_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y4_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y6_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ;
wire	\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ;
wire	\sys_resetn~combout ;
wire	\~GND~combout ;
wire	\~VCC~combout ;

wire vcc;
wire gnd;
assign vcc = 1'b1;
assign gnd = 1'b0;
wire unknown;
assign unknown = 1'bx;

alta_rio \CI_CK~input (
	.padio(CI_CK),
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\CI_CK~input_o ),
	.regout());
defparam \CI_CK~input .coord_x = 6;
defparam \CI_CK~input .coord_y = 0;
defparam \CI_CK~input .coord_z = 0;
defparam \CI_CK~input .IN_ASYNC_MODE = 1'b0;
defparam \CI_CK~input .IN_SYNC_MODE = 1'b0;
defparam \CI_CK~input .IN_POWERUP = 1'b0;
defparam \CI_CK~input .OUT_REG_MODE = 1'b0;
defparam \CI_CK~input .OUT_ASYNC_MODE = 1'b0;
defparam \CI_CK~input .OUT_SYNC_MODE = 1'b0;
defparam \CI_CK~input .OUT_POWERUP = 1'b0;
defparam \CI_CK~input .OE_REG_MODE = 1'b0;
defparam \CI_CK~input .OE_ASYNC_MODE = 1'b0;
defparam \CI_CK~input .OE_SYNC_MODE = 1'b0;
defparam \CI_CK~input .OE_POWERUP = 1'b0;
defparam \CI_CK~input .CFG_TRI_INPUT = 1'b0;
defparam \CI_CK~input .CFG_INPUT_EN = 1'b0;
defparam \CI_CK~input .CFG_PULL_UP = 1'b0;
defparam \CI_CK~input .CFG_SLR = 1'b0;
defparam \CI_CK~input .CFG_OPEN_DRAIN = 1'b0;
defparam \CI_CK~input .CFG_PDRCTRL = 4'b0100;
defparam \CI_CK~input .CFG_KEEP = 2'b00;
defparam \CI_CK~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \CI_CK~input .CFG_LVDS_SEL_CUA = 2'b00;
defparam \CI_CK~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \CI_CK~input .CFG_LVDS_IN_EN = 1'b0;
defparam \CI_CK~input .DPCLK_DELAY = 4'b0000;
defparam \CI_CK~input .OUT_DELAY = 1'b0;
defparam \CI_CK~input .IN_DATA_DELAY = 3'b000;
defparam \CI_CK~input .IN_REG_DELAY = 3'b000;

alta_rio \CI_CS~input (
	.padio(CI_CS),
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\CI_CS~input_o ),
	.regout());
defparam \CI_CS~input .coord_x = 1;
defparam \CI_CS~input .coord_y = 0;
defparam \CI_CS~input .coord_z = 3;
defparam \CI_CS~input .IN_ASYNC_MODE = 1'b0;
defparam \CI_CS~input .IN_SYNC_MODE = 1'b0;
defparam \CI_CS~input .IN_POWERUP = 1'b0;
defparam \CI_CS~input .OUT_REG_MODE = 1'b0;
defparam \CI_CS~input .OUT_ASYNC_MODE = 1'b0;
defparam \CI_CS~input .OUT_SYNC_MODE = 1'b0;
defparam \CI_CS~input .OUT_POWERUP = 1'b0;
defparam \CI_CS~input .OE_REG_MODE = 1'b0;
defparam \CI_CS~input .OE_ASYNC_MODE = 1'b0;
defparam \CI_CS~input .OE_SYNC_MODE = 1'b0;
defparam \CI_CS~input .OE_POWERUP = 1'b0;
defparam \CI_CS~input .CFG_TRI_INPUT = 1'b0;
defparam \CI_CS~input .CFG_INPUT_EN = 1'b0;
defparam \CI_CS~input .CFG_PULL_UP = 1'b0;
defparam \CI_CS~input .CFG_SLR = 1'b0;
defparam \CI_CS~input .CFG_OPEN_DRAIN = 1'b0;
defparam \CI_CS~input .CFG_PDRCTRL = 4'b0100;
defparam \CI_CS~input .CFG_KEEP = 2'b00;
defparam \CI_CS~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \CI_CS~input .CFG_LVDS_SEL_CUA = 2'b00;
defparam \CI_CS~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \CI_CS~input .CFG_LVDS_IN_EN = 1'b0;
defparam \CI_CS~input .DPCLK_DELAY = 4'b0000;
defparam \CI_CS~input .OUT_DELAY = 1'b0;
defparam \CI_CS~input .IN_DATA_DELAY = 3'b000;
defparam \CI_CS~input .IN_REG_DELAY = 3'b000;

alta_rio \CI_DAT~input (
	.padio(CI_DAT),
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\CI_DAT~input_o ),
	.regout());
defparam \CI_DAT~input .coord_x = 7;
defparam \CI_DAT~input .coord_y = 0;
defparam \CI_DAT~input .coord_z = 1;
defparam \CI_DAT~input .IN_ASYNC_MODE = 1'b0;
defparam \CI_DAT~input .IN_SYNC_MODE = 1'b0;
defparam \CI_DAT~input .IN_POWERUP = 1'b0;
defparam \CI_DAT~input .OUT_REG_MODE = 1'b0;
defparam \CI_DAT~input .OUT_ASYNC_MODE = 1'b0;
defparam \CI_DAT~input .OUT_SYNC_MODE = 1'b0;
defparam \CI_DAT~input .OUT_POWERUP = 1'b0;
defparam \CI_DAT~input .OE_REG_MODE = 1'b0;
defparam \CI_DAT~input .OE_ASYNC_MODE = 1'b0;
defparam \CI_DAT~input .OE_SYNC_MODE = 1'b0;
defparam \CI_DAT~input .OE_POWERUP = 1'b0;
defparam \CI_DAT~input .CFG_TRI_INPUT = 1'b0;
defparam \CI_DAT~input .CFG_INPUT_EN = 1'b0;
defparam \CI_DAT~input .CFG_PULL_UP = 1'b0;
defparam \CI_DAT~input .CFG_SLR = 1'b0;
defparam \CI_DAT~input .CFG_OPEN_DRAIN = 1'b0;
defparam \CI_DAT~input .CFG_PDRCTRL = 4'b0100;
defparam \CI_DAT~input .CFG_KEEP = 2'b00;
defparam \CI_DAT~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \CI_DAT~input .CFG_LVDS_SEL_CUA = 2'b00;
defparam \CI_DAT~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \CI_DAT~input .CFG_LVDS_IN_EN = 1'b0;
defparam \CI_DAT~input .DPCLK_DELAY = 4'b0000;
defparam \CI_DAT~input .OUT_DELAY = 1'b0;
defparam \CI_DAT~input .IN_DATA_DELAY = 3'b000;
defparam \CI_DAT~input .IN_REG_DELAY = 3'b000;

alta_rio \CO_CK~output (
	.padio(CO_CK),
	.datain(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \CO_CK~output .coord_x = 17;
defparam \CO_CK~output .coord_y = 0;
defparam \CO_CK~output .coord_z = 1;
defparam \CO_CK~output .IN_ASYNC_MODE = 1'b0;
defparam \CO_CK~output .IN_SYNC_MODE = 1'b0;
defparam \CO_CK~output .IN_POWERUP = 1'b0;
defparam \CO_CK~output .OUT_REG_MODE = 1'b0;
defparam \CO_CK~output .OUT_ASYNC_MODE = 1'b0;
defparam \CO_CK~output .OUT_SYNC_MODE = 1'b0;
defparam \CO_CK~output .OUT_POWERUP = 1'b0;
defparam \CO_CK~output .OE_REG_MODE = 1'b0;
defparam \CO_CK~output .OE_ASYNC_MODE = 1'b0;
defparam \CO_CK~output .OE_SYNC_MODE = 1'b0;
defparam \CO_CK~output .OE_POWERUP = 1'b0;
defparam \CO_CK~output .CFG_TRI_INPUT = 1'b0;
defparam \CO_CK~output .CFG_INPUT_EN = 1'b0;
defparam \CO_CK~output .CFG_PULL_UP = 1'b0;
defparam \CO_CK~output .CFG_SLR = 1'b0;
defparam \CO_CK~output .CFG_OPEN_DRAIN = 1'b0;
defparam \CO_CK~output .CFG_PDRCTRL = 4'b0100;
defparam \CO_CK~output .CFG_KEEP = 2'b00;
defparam \CO_CK~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \CO_CK~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \CO_CK~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \CO_CK~output .CFG_LVDS_IN_EN = 1'b0;
defparam \CO_CK~output .DPCLK_DELAY = 4'b0000;
defparam \CO_CK~output .OUT_DELAY = 1'b0;
defparam \CO_CK~output .IN_DATA_DELAY = 3'b000;
defparam \CO_CK~output .IN_REG_DELAY = 3'b000;

alta_rio \CO_CS~output (
	.padio(CO_CS),
	.datain(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \CO_CS~output .coord_x = 17;
defparam \CO_CS~output .coord_y = 0;
defparam \CO_CS~output .coord_z = 0;
defparam \CO_CS~output .IN_ASYNC_MODE = 1'b0;
defparam \CO_CS~output .IN_SYNC_MODE = 1'b0;
defparam \CO_CS~output .IN_POWERUP = 1'b0;
defparam \CO_CS~output .OUT_REG_MODE = 1'b0;
defparam \CO_CS~output .OUT_ASYNC_MODE = 1'b0;
defparam \CO_CS~output .OUT_SYNC_MODE = 1'b0;
defparam \CO_CS~output .OUT_POWERUP = 1'b0;
defparam \CO_CS~output .OE_REG_MODE = 1'b0;
defparam \CO_CS~output .OE_ASYNC_MODE = 1'b0;
defparam \CO_CS~output .OE_SYNC_MODE = 1'b0;
defparam \CO_CS~output .OE_POWERUP = 1'b0;
defparam \CO_CS~output .CFG_TRI_INPUT = 1'b0;
defparam \CO_CS~output .CFG_INPUT_EN = 1'b0;
defparam \CO_CS~output .CFG_PULL_UP = 1'b0;
defparam \CO_CS~output .CFG_SLR = 1'b0;
defparam \CO_CS~output .CFG_OPEN_DRAIN = 1'b0;
defparam \CO_CS~output .CFG_PDRCTRL = 4'b0100;
defparam \CO_CS~output .CFG_KEEP = 2'b00;
defparam \CO_CS~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \CO_CS~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \CO_CS~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \CO_CS~output .CFG_LVDS_IN_EN = 1'b0;
defparam \CO_CS~output .DPCLK_DELAY = 4'b0000;
defparam \CO_CS~output .OUT_DELAY = 1'b0;
defparam \CO_CS~output .IN_DATA_DELAY = 3'b000;
defparam \CO_CS~output .IN_REG_DELAY = 3'b000;

alta_rio \CO_DAT~output (
	.padio(CO_DAT),
	.datain(gnd),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \CO_DAT~output .coord_x = 17;
defparam \CO_DAT~output .coord_y = 0;
defparam \CO_DAT~output .coord_z = 2;
defparam \CO_DAT~output .IN_ASYNC_MODE = 1'b0;
defparam \CO_DAT~output .IN_SYNC_MODE = 1'b0;
defparam \CO_DAT~output .IN_POWERUP = 1'b0;
defparam \CO_DAT~output .OUT_REG_MODE = 1'b0;
defparam \CO_DAT~output .OUT_ASYNC_MODE = 1'b0;
defparam \CO_DAT~output .OUT_SYNC_MODE = 1'b0;
defparam \CO_DAT~output .OUT_POWERUP = 1'b0;
defparam \CO_DAT~output .OE_REG_MODE = 1'b0;
defparam \CO_DAT~output .OE_ASYNC_MODE = 1'b0;
defparam \CO_DAT~output .OE_SYNC_MODE = 1'b0;
defparam \CO_DAT~output .OE_POWERUP = 1'b0;
defparam \CO_DAT~output .CFG_TRI_INPUT = 1'b0;
defparam \CO_DAT~output .CFG_INPUT_EN = 1'b0;
defparam \CO_DAT~output .CFG_PULL_UP = 1'b0;
defparam \CO_DAT~output .CFG_SLR = 1'b0;
defparam \CO_DAT~output .CFG_OPEN_DRAIN = 1'b0;
defparam \CO_DAT~output .CFG_PDRCTRL = 4'b0100;
defparam \CO_DAT~output .CFG_KEEP = 2'b00;
defparam \CO_DAT~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \CO_DAT~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \CO_DAT~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \CO_DAT~output .CFG_LVDS_IN_EN = 1'b0;
defparam \CO_DAT~output .DPCLK_DELAY = 4'b0000;
defparam \CO_DAT~output .OUT_DELAY = 1'b0;
defparam \CO_DAT~output .IN_DATA_DELAY = 3'b000;
defparam \CO_DAT~output .IN_REG_DELAY = 3'b000;

alta_rio \D0~output (
	.padio(D0),
	.datain(\macro_inst|controller|serial|sdata_reg [0]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D0~output .coord_x = 17;
defparam \D0~output .coord_y = 13;
defparam \D0~output .coord_z = 3;
defparam \D0~output .IN_ASYNC_MODE = 1'b0;
defparam \D0~output .IN_SYNC_MODE = 1'b0;
defparam \D0~output .IN_POWERUP = 1'b0;
defparam \D0~output .OUT_REG_MODE = 1'b0;
defparam \D0~output .OUT_ASYNC_MODE = 1'b0;
defparam \D0~output .OUT_SYNC_MODE = 1'b0;
defparam \D0~output .OUT_POWERUP = 1'b0;
defparam \D0~output .OE_REG_MODE = 1'b0;
defparam \D0~output .OE_ASYNC_MODE = 1'b0;
defparam \D0~output .OE_SYNC_MODE = 1'b0;
defparam \D0~output .OE_POWERUP = 1'b0;
defparam \D0~output .CFG_TRI_INPUT = 1'b0;
defparam \D0~output .CFG_INPUT_EN = 1'b0;
defparam \D0~output .CFG_PULL_UP = 1'b0;
defparam \D0~output .CFG_SLR = 1'b0;
defparam \D0~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D0~output .CFG_PDRCTRL = 4'b0100;
defparam \D0~output .CFG_KEEP = 2'b00;
defparam \D0~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D0~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D0~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D0~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D0~output .DPCLK_DELAY = 4'b0000;
defparam \D0~output .OUT_DELAY = 1'b0;
defparam \D0~output .IN_DATA_DELAY = 3'b000;
defparam \D0~output .IN_REG_DELAY = 3'b000;

alta_rio \D10~output (
	.padio(D10),
	.datain(\macro_inst|controller|serial|sdata_reg [10]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D10~output .coord_x = 0;
defparam \D10~output .coord_y = 2;
defparam \D10~output .coord_z = 4;
defparam \D10~output .IN_ASYNC_MODE = 1'b0;
defparam \D10~output .IN_SYNC_MODE = 1'b0;
defparam \D10~output .IN_POWERUP = 1'b0;
defparam \D10~output .OUT_REG_MODE = 1'b0;
defparam \D10~output .OUT_ASYNC_MODE = 1'b0;
defparam \D10~output .OUT_SYNC_MODE = 1'b0;
defparam \D10~output .OUT_POWERUP = 1'b0;
defparam \D10~output .OE_REG_MODE = 1'b0;
defparam \D10~output .OE_ASYNC_MODE = 1'b0;
defparam \D10~output .OE_SYNC_MODE = 1'b0;
defparam \D10~output .OE_POWERUP = 1'b0;
defparam \D10~output .CFG_TRI_INPUT = 1'b0;
defparam \D10~output .CFG_INPUT_EN = 1'b0;
defparam \D10~output .CFG_PULL_UP = 1'b0;
defparam \D10~output .CFG_SLR = 1'b0;
defparam \D10~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D10~output .CFG_PDRCTRL = 4'b0100;
defparam \D10~output .CFG_KEEP = 2'b00;
defparam \D10~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D10~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D10~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D10~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D10~output .DPCLK_DELAY = 4'b0000;
defparam \D10~output .OUT_DELAY = 1'b0;
defparam \D10~output .IN_DATA_DELAY = 3'b000;
defparam \D10~output .IN_REG_DELAY = 3'b000;

alta_rio \D11~output (
	.padio(D11),
	.datain(\macro_inst|controller|serial|sdata_reg [11]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D11~output .coord_x = 0;
defparam \D11~output .coord_y = 2;
defparam \D11~output .coord_z = 5;
defparam \D11~output .IN_ASYNC_MODE = 1'b0;
defparam \D11~output .IN_SYNC_MODE = 1'b0;
defparam \D11~output .IN_POWERUP = 1'b0;
defparam \D11~output .OUT_REG_MODE = 1'b0;
defparam \D11~output .OUT_ASYNC_MODE = 1'b0;
defparam \D11~output .OUT_SYNC_MODE = 1'b0;
defparam \D11~output .OUT_POWERUP = 1'b0;
defparam \D11~output .OE_REG_MODE = 1'b0;
defparam \D11~output .OE_ASYNC_MODE = 1'b0;
defparam \D11~output .OE_SYNC_MODE = 1'b0;
defparam \D11~output .OE_POWERUP = 1'b0;
defparam \D11~output .CFG_TRI_INPUT = 1'b0;
defparam \D11~output .CFG_INPUT_EN = 1'b0;
defparam \D11~output .CFG_PULL_UP = 1'b0;
defparam \D11~output .CFG_SLR = 1'b0;
defparam \D11~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D11~output .CFG_PDRCTRL = 4'b0100;
defparam \D11~output .CFG_KEEP = 2'b00;
defparam \D11~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D11~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D11~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D11~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D11~output .DPCLK_DELAY = 4'b0000;
defparam \D11~output .OUT_DELAY = 1'b0;
defparam \D11~output .IN_DATA_DELAY = 3'b000;
defparam \D11~output .IN_REG_DELAY = 3'b000;

alta_rio \D12~output (
	.padio(D12),
	.datain(\macro_inst|controller|serial|sdata_reg [12]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D12~output .coord_x = 18;
defparam \D12~output .coord_y = 0;
defparam \D12~output .coord_z = 0;
defparam \D12~output .IN_ASYNC_MODE = 1'b0;
defparam \D12~output .IN_SYNC_MODE = 1'b0;
defparam \D12~output .IN_POWERUP = 1'b0;
defparam \D12~output .OUT_REG_MODE = 1'b0;
defparam \D12~output .OUT_ASYNC_MODE = 1'b0;
defparam \D12~output .OUT_SYNC_MODE = 1'b0;
defparam \D12~output .OUT_POWERUP = 1'b0;
defparam \D12~output .OE_REG_MODE = 1'b0;
defparam \D12~output .OE_ASYNC_MODE = 1'b0;
defparam \D12~output .OE_SYNC_MODE = 1'b0;
defparam \D12~output .OE_POWERUP = 1'b0;
defparam \D12~output .CFG_TRI_INPUT = 1'b0;
defparam \D12~output .CFG_INPUT_EN = 1'b0;
defparam \D12~output .CFG_PULL_UP = 1'b0;
defparam \D12~output .CFG_SLR = 1'b0;
defparam \D12~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D12~output .CFG_PDRCTRL = 4'b0100;
defparam \D12~output .CFG_KEEP = 2'b00;
defparam \D12~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D12~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D12~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D12~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D12~output .DPCLK_DELAY = 4'b0000;
defparam \D12~output .OUT_DELAY = 1'b0;
defparam \D12~output .IN_DATA_DELAY = 3'b000;
defparam \D12~output .IN_REG_DELAY = 3'b000;

alta_rio \D13~output (
	.padio(D13),
	.datain(\macro_inst|controller|serial|sdata_reg [13]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D13~output .coord_x = 18;
defparam \D13~output .coord_y = 0;
defparam \D13~output .coord_z = 1;
defparam \D13~output .IN_ASYNC_MODE = 1'b0;
defparam \D13~output .IN_SYNC_MODE = 1'b0;
defparam \D13~output .IN_POWERUP = 1'b0;
defparam \D13~output .OUT_REG_MODE = 1'b0;
defparam \D13~output .OUT_ASYNC_MODE = 1'b0;
defparam \D13~output .OUT_SYNC_MODE = 1'b0;
defparam \D13~output .OUT_POWERUP = 1'b0;
defparam \D13~output .OE_REG_MODE = 1'b0;
defparam \D13~output .OE_ASYNC_MODE = 1'b0;
defparam \D13~output .OE_SYNC_MODE = 1'b0;
defparam \D13~output .OE_POWERUP = 1'b0;
defparam \D13~output .CFG_TRI_INPUT = 1'b0;
defparam \D13~output .CFG_INPUT_EN = 1'b0;
defparam \D13~output .CFG_PULL_UP = 1'b0;
defparam \D13~output .CFG_SLR = 1'b0;
defparam \D13~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D13~output .CFG_PDRCTRL = 4'b0100;
defparam \D13~output .CFG_KEEP = 2'b00;
defparam \D13~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D13~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D13~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D13~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D13~output .DPCLK_DELAY = 4'b0000;
defparam \D13~output .OUT_DELAY = 1'b0;
defparam \D13~output .IN_DATA_DELAY = 3'b000;
defparam \D13~output .IN_REG_DELAY = 3'b000;

alta_rio \D14~output (
	.padio(D14),
	.datain(\macro_inst|controller|serial|sdata_reg [14]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D14~output .coord_x = 18;
defparam \D14~output .coord_y = 13;
defparam \D14~output .coord_z = 2;
defparam \D14~output .IN_ASYNC_MODE = 1'b0;
defparam \D14~output .IN_SYNC_MODE = 1'b0;
defparam \D14~output .IN_POWERUP = 1'b0;
defparam \D14~output .OUT_REG_MODE = 1'b0;
defparam \D14~output .OUT_ASYNC_MODE = 1'b0;
defparam \D14~output .OUT_SYNC_MODE = 1'b0;
defparam \D14~output .OUT_POWERUP = 1'b0;
defparam \D14~output .OE_REG_MODE = 1'b0;
defparam \D14~output .OE_ASYNC_MODE = 1'b0;
defparam \D14~output .OE_SYNC_MODE = 1'b0;
defparam \D14~output .OE_POWERUP = 1'b0;
defparam \D14~output .CFG_TRI_INPUT = 1'b0;
defparam \D14~output .CFG_INPUT_EN = 1'b0;
defparam \D14~output .CFG_PULL_UP = 1'b0;
defparam \D14~output .CFG_SLR = 1'b0;
defparam \D14~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D14~output .CFG_PDRCTRL = 4'b0100;
defparam \D14~output .CFG_KEEP = 2'b00;
defparam \D14~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D14~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D14~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D14~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D14~output .DPCLK_DELAY = 4'b0000;
defparam \D14~output .OUT_DELAY = 1'b0;
defparam \D14~output .IN_DATA_DELAY = 3'b000;
defparam \D14~output .IN_REG_DELAY = 3'b000;

alta_rio \D15~output (
	.padio(D15),
	.datain(\macro_inst|controller|serial|sdata_reg [15]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D15~output .coord_x = 18;
defparam \D15~output .coord_y = 13;
defparam \D15~output .coord_z = 1;
defparam \D15~output .IN_ASYNC_MODE = 1'b0;
defparam \D15~output .IN_SYNC_MODE = 1'b0;
defparam \D15~output .IN_POWERUP = 1'b0;
defparam \D15~output .OUT_REG_MODE = 1'b0;
defparam \D15~output .OUT_ASYNC_MODE = 1'b0;
defparam \D15~output .OUT_SYNC_MODE = 1'b0;
defparam \D15~output .OUT_POWERUP = 1'b0;
defparam \D15~output .OE_REG_MODE = 1'b0;
defparam \D15~output .OE_ASYNC_MODE = 1'b0;
defparam \D15~output .OE_SYNC_MODE = 1'b0;
defparam \D15~output .OE_POWERUP = 1'b0;
defparam \D15~output .CFG_TRI_INPUT = 1'b0;
defparam \D15~output .CFG_INPUT_EN = 1'b0;
defparam \D15~output .CFG_PULL_UP = 1'b0;
defparam \D15~output .CFG_SLR = 1'b0;
defparam \D15~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D15~output .CFG_PDRCTRL = 4'b0100;
defparam \D15~output .CFG_KEEP = 2'b00;
defparam \D15~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D15~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D15~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D15~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D15~output .DPCLK_DELAY = 4'b0000;
defparam \D15~output .OUT_DELAY = 1'b0;
defparam \D15~output .IN_DATA_DELAY = 3'b000;
defparam \D15~output .IN_REG_DELAY = 3'b000;

alta_rio \D16~output (
	.padio(D16),
	.datain(\macro_inst|controller|serial|sdata_reg [16]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D16~output .coord_x = 19;
defparam \D16~output .coord_y = 0;
defparam \D16~output .coord_z = 3;
defparam \D16~output .IN_ASYNC_MODE = 1'b0;
defparam \D16~output .IN_SYNC_MODE = 1'b0;
defparam \D16~output .IN_POWERUP = 1'b0;
defparam \D16~output .OUT_REG_MODE = 1'b0;
defparam \D16~output .OUT_ASYNC_MODE = 1'b0;
defparam \D16~output .OUT_SYNC_MODE = 1'b0;
defparam \D16~output .OUT_POWERUP = 1'b0;
defparam \D16~output .OE_REG_MODE = 1'b0;
defparam \D16~output .OE_ASYNC_MODE = 1'b0;
defparam \D16~output .OE_SYNC_MODE = 1'b0;
defparam \D16~output .OE_POWERUP = 1'b0;
defparam \D16~output .CFG_TRI_INPUT = 1'b0;
defparam \D16~output .CFG_INPUT_EN = 1'b0;
defparam \D16~output .CFG_PULL_UP = 1'b0;
defparam \D16~output .CFG_SLR = 1'b0;
defparam \D16~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D16~output .CFG_PDRCTRL = 4'b0100;
defparam \D16~output .CFG_KEEP = 2'b00;
defparam \D16~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D16~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D16~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D16~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D16~output .DPCLK_DELAY = 4'b0000;
defparam \D16~output .OUT_DELAY = 1'b0;
defparam \D16~output .IN_DATA_DELAY = 3'b000;
defparam \D16~output .IN_REG_DELAY = 3'b000;

alta_rio \D17~output (
	.padio(D17),
	.datain(\macro_inst|controller|serial|sdata_reg [17]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D17~output .coord_x = 22;
defparam \D17~output .coord_y = 2;
defparam \D17~output .coord_z = 3;
defparam \D17~output .IN_ASYNC_MODE = 1'b0;
defparam \D17~output .IN_SYNC_MODE = 1'b0;
defparam \D17~output .IN_POWERUP = 1'b0;
defparam \D17~output .OUT_REG_MODE = 1'b0;
defparam \D17~output .OUT_ASYNC_MODE = 1'b0;
defparam \D17~output .OUT_SYNC_MODE = 1'b0;
defparam \D17~output .OUT_POWERUP = 1'b0;
defparam \D17~output .OE_REG_MODE = 1'b0;
defparam \D17~output .OE_ASYNC_MODE = 1'b0;
defparam \D17~output .OE_SYNC_MODE = 1'b0;
defparam \D17~output .OE_POWERUP = 1'b0;
defparam \D17~output .CFG_TRI_INPUT = 1'b0;
defparam \D17~output .CFG_INPUT_EN = 1'b0;
defparam \D17~output .CFG_PULL_UP = 1'b0;
defparam \D17~output .CFG_SLR = 1'b0;
defparam \D17~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D17~output .CFG_PDRCTRL = 4'b0100;
defparam \D17~output .CFG_KEEP = 2'b00;
defparam \D17~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D17~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D17~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D17~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D17~output .DPCLK_DELAY = 4'b0000;
defparam \D17~output .OUT_DELAY = 1'b0;
defparam \D17~output .IN_DATA_DELAY = 3'b000;
defparam \D17~output .IN_REG_DELAY = 3'b000;

alta_rio \D18~output (
	.padio(D18),
	.datain(\macro_inst|controller|serial|sdata_reg [18]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D18~output .coord_x = 19;
defparam \D18~output .coord_y = 13;
defparam \D18~output .coord_z = 1;
defparam \D18~output .IN_ASYNC_MODE = 1'b0;
defparam \D18~output .IN_SYNC_MODE = 1'b0;
defparam \D18~output .IN_POWERUP = 1'b0;
defparam \D18~output .OUT_REG_MODE = 1'b0;
defparam \D18~output .OUT_ASYNC_MODE = 1'b0;
defparam \D18~output .OUT_SYNC_MODE = 1'b0;
defparam \D18~output .OUT_POWERUP = 1'b0;
defparam \D18~output .OE_REG_MODE = 1'b0;
defparam \D18~output .OE_ASYNC_MODE = 1'b0;
defparam \D18~output .OE_SYNC_MODE = 1'b0;
defparam \D18~output .OE_POWERUP = 1'b0;
defparam \D18~output .CFG_TRI_INPUT = 1'b0;
defparam \D18~output .CFG_INPUT_EN = 1'b0;
defparam \D18~output .CFG_PULL_UP = 1'b0;
defparam \D18~output .CFG_SLR = 1'b0;
defparam \D18~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D18~output .CFG_PDRCTRL = 4'b0100;
defparam \D18~output .CFG_KEEP = 2'b00;
defparam \D18~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D18~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D18~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D18~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D18~output .DPCLK_DELAY = 4'b0000;
defparam \D18~output .OUT_DELAY = 1'b0;
defparam \D18~output .IN_DATA_DELAY = 3'b000;
defparam \D18~output .IN_REG_DELAY = 3'b000;

alta_rio \D19~output (
	.padio(D19),
	.datain(\macro_inst|controller|serial|sdata_reg [19]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D19~output .coord_x = 19;
defparam \D19~output .coord_y = 13;
defparam \D19~output .coord_z = 0;
defparam \D19~output .IN_ASYNC_MODE = 1'b0;
defparam \D19~output .IN_SYNC_MODE = 1'b0;
defparam \D19~output .IN_POWERUP = 1'b0;
defparam \D19~output .OUT_REG_MODE = 1'b0;
defparam \D19~output .OUT_ASYNC_MODE = 1'b0;
defparam \D19~output .OUT_SYNC_MODE = 1'b0;
defparam \D19~output .OUT_POWERUP = 1'b0;
defparam \D19~output .OE_REG_MODE = 1'b0;
defparam \D19~output .OE_ASYNC_MODE = 1'b0;
defparam \D19~output .OE_SYNC_MODE = 1'b0;
defparam \D19~output .OE_POWERUP = 1'b0;
defparam \D19~output .CFG_TRI_INPUT = 1'b0;
defparam \D19~output .CFG_INPUT_EN = 1'b0;
defparam \D19~output .CFG_PULL_UP = 1'b0;
defparam \D19~output .CFG_SLR = 1'b0;
defparam \D19~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D19~output .CFG_PDRCTRL = 4'b0100;
defparam \D19~output .CFG_KEEP = 2'b00;
defparam \D19~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D19~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D19~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D19~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D19~output .DPCLK_DELAY = 4'b0000;
defparam \D19~output .OUT_DELAY = 1'b0;
defparam \D19~output .IN_DATA_DELAY = 3'b000;
defparam \D19~output .IN_REG_DELAY = 3'b000;

alta_rio \D1~output (
	.padio(D1),
	.datain(\macro_inst|controller|serial|sdata_reg [1]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D1~output .coord_x = 17;
defparam \D1~output .coord_y = 13;
defparam \D1~output .coord_z = 2;
defparam \D1~output .IN_ASYNC_MODE = 1'b0;
defparam \D1~output .IN_SYNC_MODE = 1'b0;
defparam \D1~output .IN_POWERUP = 1'b0;
defparam \D1~output .OUT_REG_MODE = 1'b0;
defparam \D1~output .OUT_ASYNC_MODE = 1'b0;
defparam \D1~output .OUT_SYNC_MODE = 1'b0;
defparam \D1~output .OUT_POWERUP = 1'b0;
defparam \D1~output .OE_REG_MODE = 1'b0;
defparam \D1~output .OE_ASYNC_MODE = 1'b0;
defparam \D1~output .OE_SYNC_MODE = 1'b0;
defparam \D1~output .OE_POWERUP = 1'b0;
defparam \D1~output .CFG_TRI_INPUT = 1'b0;
defparam \D1~output .CFG_INPUT_EN = 1'b0;
defparam \D1~output .CFG_PULL_UP = 1'b0;
defparam \D1~output .CFG_SLR = 1'b0;
defparam \D1~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D1~output .CFG_PDRCTRL = 4'b0100;
defparam \D1~output .CFG_KEEP = 2'b00;
defparam \D1~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D1~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D1~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D1~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D1~output .DPCLK_DELAY = 4'b0000;
defparam \D1~output .OUT_DELAY = 1'b0;
defparam \D1~output .IN_DATA_DELAY = 3'b000;
defparam \D1~output .IN_REG_DELAY = 3'b000;

alta_rio \D20~output (
	.padio(D20),
	.datain(\macro_inst|controller|serial|sdata_reg [20]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D20~output .coord_x = 22;
defparam \D20~output .coord_y = 3;
defparam \D20~output .coord_z = 2;
defparam \D20~output .IN_ASYNC_MODE = 1'b0;
defparam \D20~output .IN_SYNC_MODE = 1'b0;
defparam \D20~output .IN_POWERUP = 1'b0;
defparam \D20~output .OUT_REG_MODE = 1'b0;
defparam \D20~output .OUT_ASYNC_MODE = 1'b0;
defparam \D20~output .OUT_SYNC_MODE = 1'b0;
defparam \D20~output .OUT_POWERUP = 1'b0;
defparam \D20~output .OE_REG_MODE = 1'b0;
defparam \D20~output .OE_ASYNC_MODE = 1'b0;
defparam \D20~output .OE_SYNC_MODE = 1'b0;
defparam \D20~output .OE_POWERUP = 1'b0;
defparam \D20~output .CFG_TRI_INPUT = 1'b0;
defparam \D20~output .CFG_INPUT_EN = 1'b0;
defparam \D20~output .CFG_PULL_UP = 1'b0;
defparam \D20~output .CFG_SLR = 1'b0;
defparam \D20~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D20~output .CFG_PDRCTRL = 4'b0100;
defparam \D20~output .CFG_KEEP = 2'b00;
defparam \D20~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D20~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D20~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D20~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D20~output .DPCLK_DELAY = 4'b0000;
defparam \D20~output .OUT_DELAY = 1'b0;
defparam \D20~output .IN_DATA_DELAY = 3'b000;
defparam \D20~output .IN_REG_DELAY = 3'b000;

alta_rio \D21~output (
	.padio(D21),
	.datain(\macro_inst|controller|serial|sdata_reg [21]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D21~output .coord_x = 22;
defparam \D21~output .coord_y = 3;
defparam \D21~output .coord_z = 1;
defparam \D21~output .IN_ASYNC_MODE = 1'b0;
defparam \D21~output .IN_SYNC_MODE = 1'b0;
defparam \D21~output .IN_POWERUP = 1'b0;
defparam \D21~output .OUT_REG_MODE = 1'b0;
defparam \D21~output .OUT_ASYNC_MODE = 1'b0;
defparam \D21~output .OUT_SYNC_MODE = 1'b0;
defparam \D21~output .OUT_POWERUP = 1'b0;
defparam \D21~output .OE_REG_MODE = 1'b0;
defparam \D21~output .OE_ASYNC_MODE = 1'b0;
defparam \D21~output .OE_SYNC_MODE = 1'b0;
defparam \D21~output .OE_POWERUP = 1'b0;
defparam \D21~output .CFG_TRI_INPUT = 1'b0;
defparam \D21~output .CFG_INPUT_EN = 1'b0;
defparam \D21~output .CFG_PULL_UP = 1'b0;
defparam \D21~output .CFG_SLR = 1'b0;
defparam \D21~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D21~output .CFG_PDRCTRL = 4'b0100;
defparam \D21~output .CFG_KEEP = 2'b00;
defparam \D21~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D21~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D21~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D21~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D21~output .DPCLK_DELAY = 4'b0000;
defparam \D21~output .OUT_DELAY = 1'b0;
defparam \D21~output .IN_DATA_DELAY = 3'b000;
defparam \D21~output .IN_REG_DELAY = 3'b000;

alta_rio \D22~output (
	.padio(D22),
	.datain(\macro_inst|controller|serial|sdata_reg [22]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D22~output .coord_x = 20;
defparam \D22~output .coord_y = 13;
defparam \D22~output .coord_z = 3;
defparam \D22~output .IN_ASYNC_MODE = 1'b0;
defparam \D22~output .IN_SYNC_MODE = 1'b0;
defparam \D22~output .IN_POWERUP = 1'b0;
defparam \D22~output .OUT_REG_MODE = 1'b0;
defparam \D22~output .OUT_ASYNC_MODE = 1'b0;
defparam \D22~output .OUT_SYNC_MODE = 1'b0;
defparam \D22~output .OUT_POWERUP = 1'b0;
defparam \D22~output .OE_REG_MODE = 1'b0;
defparam \D22~output .OE_ASYNC_MODE = 1'b0;
defparam \D22~output .OE_SYNC_MODE = 1'b0;
defparam \D22~output .OE_POWERUP = 1'b0;
defparam \D22~output .CFG_TRI_INPUT = 1'b0;
defparam \D22~output .CFG_INPUT_EN = 1'b0;
defparam \D22~output .CFG_PULL_UP = 1'b0;
defparam \D22~output .CFG_SLR = 1'b0;
defparam \D22~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D22~output .CFG_PDRCTRL = 4'b0100;
defparam \D22~output .CFG_KEEP = 2'b00;
defparam \D22~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D22~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D22~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D22~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D22~output .DPCLK_DELAY = 4'b0000;
defparam \D22~output .OUT_DELAY = 1'b0;
defparam \D22~output .IN_DATA_DELAY = 3'b000;
defparam \D22~output .IN_REG_DELAY = 3'b000;

alta_rio \D23~output (
	.padio(D23),
	.datain(\macro_inst|controller|serial|sdata_reg [23]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D23~output .coord_x = 19;
defparam \D23~output .coord_y = 13;
defparam \D23~output .coord_z = 3;
defparam \D23~output .IN_ASYNC_MODE = 1'b0;
defparam \D23~output .IN_SYNC_MODE = 1'b0;
defparam \D23~output .IN_POWERUP = 1'b0;
defparam \D23~output .OUT_REG_MODE = 1'b0;
defparam \D23~output .OUT_ASYNC_MODE = 1'b0;
defparam \D23~output .OUT_SYNC_MODE = 1'b0;
defparam \D23~output .OUT_POWERUP = 1'b0;
defparam \D23~output .OE_REG_MODE = 1'b0;
defparam \D23~output .OE_ASYNC_MODE = 1'b0;
defparam \D23~output .OE_SYNC_MODE = 1'b0;
defparam \D23~output .OE_POWERUP = 1'b0;
defparam \D23~output .CFG_TRI_INPUT = 1'b0;
defparam \D23~output .CFG_INPUT_EN = 1'b0;
defparam \D23~output .CFG_PULL_UP = 1'b0;
defparam \D23~output .CFG_SLR = 1'b0;
defparam \D23~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D23~output .CFG_PDRCTRL = 4'b0100;
defparam \D23~output .CFG_KEEP = 2'b00;
defparam \D23~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D23~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D23~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D23~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D23~output .DPCLK_DELAY = 4'b0000;
defparam \D23~output .OUT_DELAY = 1'b0;
defparam \D23~output .IN_DATA_DELAY = 3'b000;
defparam \D23~output .IN_REG_DELAY = 3'b000;

alta_rio \D2~output (
	.padio(D2),
	.datain(\macro_inst|controller|serial|sdata_reg [2]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D2~output .coord_x = 1;
defparam \D2~output .coord_y = 0;
defparam \D2~output .coord_z = 1;
defparam \D2~output .IN_ASYNC_MODE = 1'b0;
defparam \D2~output .IN_SYNC_MODE = 1'b0;
defparam \D2~output .IN_POWERUP = 1'b0;
defparam \D2~output .OUT_REG_MODE = 1'b0;
defparam \D2~output .OUT_ASYNC_MODE = 1'b0;
defparam \D2~output .OUT_SYNC_MODE = 1'b0;
defparam \D2~output .OUT_POWERUP = 1'b0;
defparam \D2~output .OE_REG_MODE = 1'b0;
defparam \D2~output .OE_ASYNC_MODE = 1'b0;
defparam \D2~output .OE_SYNC_MODE = 1'b0;
defparam \D2~output .OE_POWERUP = 1'b0;
defparam \D2~output .CFG_TRI_INPUT = 1'b0;
defparam \D2~output .CFG_INPUT_EN = 1'b0;
defparam \D2~output .CFG_PULL_UP = 1'b0;
defparam \D2~output .CFG_SLR = 1'b0;
defparam \D2~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D2~output .CFG_PDRCTRL = 4'b0100;
defparam \D2~output .CFG_KEEP = 2'b00;
defparam \D2~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D2~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D2~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D2~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D2~output .DPCLK_DELAY = 4'b0000;
defparam \D2~output .OUT_DELAY = 1'b0;
defparam \D2~output .IN_DATA_DELAY = 3'b000;
defparam \D2~output .IN_REG_DELAY = 3'b000;

alta_rio \D3~output (
	.padio(D3),
	.datain(\macro_inst|controller|serial|sdata_reg [3]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D3~output .coord_x = 1;
defparam \D3~output .coord_y = 0;
defparam \D3~output .coord_z = 2;
defparam \D3~output .IN_ASYNC_MODE = 1'b0;
defparam \D3~output .IN_SYNC_MODE = 1'b0;
defparam \D3~output .IN_POWERUP = 1'b0;
defparam \D3~output .OUT_REG_MODE = 1'b0;
defparam \D3~output .OUT_ASYNC_MODE = 1'b0;
defparam \D3~output .OUT_SYNC_MODE = 1'b0;
defparam \D3~output .OUT_POWERUP = 1'b0;
defparam \D3~output .OE_REG_MODE = 1'b0;
defparam \D3~output .OE_ASYNC_MODE = 1'b0;
defparam \D3~output .OE_SYNC_MODE = 1'b0;
defparam \D3~output .OE_POWERUP = 1'b0;
defparam \D3~output .CFG_TRI_INPUT = 1'b0;
defparam \D3~output .CFG_INPUT_EN = 1'b0;
defparam \D3~output .CFG_PULL_UP = 1'b0;
defparam \D3~output .CFG_SLR = 1'b0;
defparam \D3~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D3~output .CFG_PDRCTRL = 4'b0100;
defparam \D3~output .CFG_KEEP = 2'b00;
defparam \D3~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D3~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D3~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D3~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D3~output .DPCLK_DELAY = 4'b0000;
defparam \D3~output .OUT_DELAY = 1'b0;
defparam \D3~output .IN_DATA_DELAY = 3'b000;
defparam \D3~output .IN_REG_DELAY = 3'b000;

alta_rio \D4~output (
	.padio(D4),
	.datain(\macro_inst|controller|serial|sdata_reg [4]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D4~output .coord_x = 16;
defparam \D4~output .coord_y = 13;
defparam \D4~output .coord_z = 1;
defparam \D4~output .IN_ASYNC_MODE = 1'b0;
defparam \D4~output .IN_SYNC_MODE = 1'b0;
defparam \D4~output .IN_POWERUP = 1'b0;
defparam \D4~output .OUT_REG_MODE = 1'b0;
defparam \D4~output .OUT_ASYNC_MODE = 1'b0;
defparam \D4~output .OUT_SYNC_MODE = 1'b0;
defparam \D4~output .OUT_POWERUP = 1'b0;
defparam \D4~output .OE_REG_MODE = 1'b0;
defparam \D4~output .OE_ASYNC_MODE = 1'b0;
defparam \D4~output .OE_SYNC_MODE = 1'b0;
defparam \D4~output .OE_POWERUP = 1'b0;
defparam \D4~output .CFG_TRI_INPUT = 1'b0;
defparam \D4~output .CFG_INPUT_EN = 1'b0;
defparam \D4~output .CFG_PULL_UP = 1'b0;
defparam \D4~output .CFG_SLR = 1'b0;
defparam \D4~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D4~output .CFG_PDRCTRL = 4'b0100;
defparam \D4~output .CFG_KEEP = 2'b00;
defparam \D4~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D4~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D4~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D4~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D4~output .DPCLK_DELAY = 4'b0000;
defparam \D4~output .OUT_DELAY = 1'b0;
defparam \D4~output .IN_DATA_DELAY = 3'b000;
defparam \D4~output .IN_REG_DELAY = 3'b000;

alta_rio \D5~output (
	.padio(D5),
	.datain(\macro_inst|controller|serial|sdata_reg [5]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D5~output .coord_x = 14;
defparam \D5~output .coord_y = 13;
defparam \D5~output .coord_z = 0;
defparam \D5~output .IN_ASYNC_MODE = 1'b0;
defparam \D5~output .IN_SYNC_MODE = 1'b0;
defparam \D5~output .IN_POWERUP = 1'b0;
defparam \D5~output .OUT_REG_MODE = 1'b0;
defparam \D5~output .OUT_ASYNC_MODE = 1'b0;
defparam \D5~output .OUT_SYNC_MODE = 1'b0;
defparam \D5~output .OUT_POWERUP = 1'b0;
defparam \D5~output .OE_REG_MODE = 1'b0;
defparam \D5~output .OE_ASYNC_MODE = 1'b0;
defparam \D5~output .OE_SYNC_MODE = 1'b0;
defparam \D5~output .OE_POWERUP = 1'b0;
defparam \D5~output .CFG_TRI_INPUT = 1'b0;
defparam \D5~output .CFG_INPUT_EN = 1'b0;
defparam \D5~output .CFG_PULL_UP = 1'b0;
defparam \D5~output .CFG_SLR = 1'b0;
defparam \D5~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D5~output .CFG_PDRCTRL = 4'b0100;
defparam \D5~output .CFG_KEEP = 2'b00;
defparam \D5~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D5~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D5~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D5~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D5~output .DPCLK_DELAY = 4'b0000;
defparam \D5~output .OUT_DELAY = 1'b0;
defparam \D5~output .IN_DATA_DELAY = 3'b000;
defparam \D5~output .IN_REG_DELAY = 3'b000;

alta_rio \D6~output (
	.padio(D6),
	.datain(\macro_inst|controller|serial|sdata_reg [6]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D6~output .coord_x = 0;
defparam \D6~output .coord_y = 1;
defparam \D6~output .coord_z = 2;
defparam \D6~output .IN_ASYNC_MODE = 1'b0;
defparam \D6~output .IN_SYNC_MODE = 1'b0;
defparam \D6~output .IN_POWERUP = 1'b0;
defparam \D6~output .OUT_REG_MODE = 1'b0;
defparam \D6~output .OUT_ASYNC_MODE = 1'b0;
defparam \D6~output .OUT_SYNC_MODE = 1'b0;
defparam \D6~output .OUT_POWERUP = 1'b0;
defparam \D6~output .OE_REG_MODE = 1'b0;
defparam \D6~output .OE_ASYNC_MODE = 1'b0;
defparam \D6~output .OE_SYNC_MODE = 1'b0;
defparam \D6~output .OE_POWERUP = 1'b0;
defparam \D6~output .CFG_TRI_INPUT = 1'b0;
defparam \D6~output .CFG_INPUT_EN = 1'b0;
defparam \D6~output .CFG_PULL_UP = 1'b0;
defparam \D6~output .CFG_SLR = 1'b0;
defparam \D6~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D6~output .CFG_PDRCTRL = 4'b0100;
defparam \D6~output .CFG_KEEP = 2'b00;
defparam \D6~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D6~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D6~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D6~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D6~output .DPCLK_DELAY = 4'b0000;
defparam \D6~output .OUT_DELAY = 1'b0;
defparam \D6~output .IN_DATA_DELAY = 3'b000;
defparam \D6~output .IN_REG_DELAY = 3'b000;

alta_rio \D7~output (
	.padio(D7),
	.datain(\macro_inst|controller|serial|sdata_reg [7]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D7~output .coord_x = 0;
defparam \D7~output .coord_y = 1;
defparam \D7~output .coord_z = 3;
defparam \D7~output .IN_ASYNC_MODE = 1'b0;
defparam \D7~output .IN_SYNC_MODE = 1'b0;
defparam \D7~output .IN_POWERUP = 1'b0;
defparam \D7~output .OUT_REG_MODE = 1'b0;
defparam \D7~output .OUT_ASYNC_MODE = 1'b0;
defparam \D7~output .OUT_SYNC_MODE = 1'b0;
defparam \D7~output .OUT_POWERUP = 1'b0;
defparam \D7~output .OE_REG_MODE = 1'b0;
defparam \D7~output .OE_ASYNC_MODE = 1'b0;
defparam \D7~output .OE_SYNC_MODE = 1'b0;
defparam \D7~output .OE_POWERUP = 1'b0;
defparam \D7~output .CFG_TRI_INPUT = 1'b0;
defparam \D7~output .CFG_INPUT_EN = 1'b0;
defparam \D7~output .CFG_PULL_UP = 1'b0;
defparam \D7~output .CFG_SLR = 1'b0;
defparam \D7~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D7~output .CFG_PDRCTRL = 4'b0100;
defparam \D7~output .CFG_KEEP = 2'b00;
defparam \D7~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D7~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D7~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D7~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D7~output .DPCLK_DELAY = 4'b0000;
defparam \D7~output .OUT_DELAY = 1'b0;
defparam \D7~output .IN_DATA_DELAY = 3'b000;
defparam \D7~output .IN_REG_DELAY = 3'b000;

alta_rio \D8~output (
	.padio(D8),
	.datain(\macro_inst|controller|serial|sdata_reg [8]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D8~output .coord_x = 0;
defparam \D8~output .coord_y = 4;
defparam \D8~output .coord_z = 1;
defparam \D8~output .IN_ASYNC_MODE = 1'b0;
defparam \D8~output .IN_SYNC_MODE = 1'b0;
defparam \D8~output .IN_POWERUP = 1'b0;
defparam \D8~output .OUT_REG_MODE = 1'b0;
defparam \D8~output .OUT_ASYNC_MODE = 1'b0;
defparam \D8~output .OUT_SYNC_MODE = 1'b0;
defparam \D8~output .OUT_POWERUP = 1'b0;
defparam \D8~output .OE_REG_MODE = 1'b0;
defparam \D8~output .OE_ASYNC_MODE = 1'b0;
defparam \D8~output .OE_SYNC_MODE = 1'b0;
defparam \D8~output .OE_POWERUP = 1'b0;
defparam \D8~output .CFG_TRI_INPUT = 1'b0;
defparam \D8~output .CFG_INPUT_EN = 1'b0;
defparam \D8~output .CFG_PULL_UP = 1'b0;
defparam \D8~output .CFG_SLR = 1'b0;
defparam \D8~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D8~output .CFG_PDRCTRL = 4'b0100;
defparam \D8~output .CFG_KEEP = 2'b00;
defparam \D8~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D8~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D8~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D8~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D8~output .DPCLK_DELAY = 4'b0000;
defparam \D8~output .OUT_DELAY = 1'b0;
defparam \D8~output .IN_DATA_DELAY = 3'b000;
defparam \D8~output .IN_REG_DELAY = 3'b000;

alta_rio \D9~output (
	.padio(D9),
	.datain(\macro_inst|controller|serial|sdata_reg [9]),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \D9~output .coord_x = 0;
defparam \D9~output .coord_y = 4;
defparam \D9~output .coord_z = 2;
defparam \D9~output .IN_ASYNC_MODE = 1'b0;
defparam \D9~output .IN_SYNC_MODE = 1'b0;
defparam \D9~output .IN_POWERUP = 1'b0;
defparam \D9~output .OUT_REG_MODE = 1'b0;
defparam \D9~output .OUT_ASYNC_MODE = 1'b0;
defparam \D9~output .OUT_SYNC_MODE = 1'b0;
defparam \D9~output .OUT_POWERUP = 1'b0;
defparam \D9~output .OE_REG_MODE = 1'b0;
defparam \D9~output .OE_ASYNC_MODE = 1'b0;
defparam \D9~output .OE_SYNC_MODE = 1'b0;
defparam \D9~output .OE_POWERUP = 1'b0;
defparam \D9~output .CFG_TRI_INPUT = 1'b0;
defparam \D9~output .CFG_INPUT_EN = 1'b0;
defparam \D9~output .CFG_PULL_UP = 1'b0;
defparam \D9~output .CFG_SLR = 1'b0;
defparam \D9~output .CFG_OPEN_DRAIN = 1'b0;
defparam \D9~output .CFG_PDRCTRL = 4'b0100;
defparam \D9~output .CFG_KEEP = 2'b00;
defparam \D9~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \D9~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \D9~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \D9~output .CFG_LVDS_IN_EN = 1'b0;
defparam \D9~output .DPCLK_DELAY = 4'b0000;
defparam \D9~output .OUT_DELAY = 1'b0;
defparam \D9~output .IN_DATA_DELAY = 3'b000;
defparam \D9~output .IN_REG_DELAY = 3'b000;

alta_rio \LM_CK~output (
	.padio(LM_CK),
	.datain(\macro_inst|serial_lim_input_inst|shift~combout ),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \LM_CK~output .coord_x = 0;
defparam \LM_CK~output .coord_y = 2;
defparam \LM_CK~output .coord_z = 1;
defparam \LM_CK~output .IN_ASYNC_MODE = 1'b0;
defparam \LM_CK~output .IN_SYNC_MODE = 1'b0;
defparam \LM_CK~output .IN_POWERUP = 1'b0;
defparam \LM_CK~output .OUT_REG_MODE = 1'b0;
defparam \LM_CK~output .OUT_ASYNC_MODE = 1'b0;
defparam \LM_CK~output .OUT_SYNC_MODE = 1'b0;
defparam \LM_CK~output .OUT_POWERUP = 1'b0;
defparam \LM_CK~output .OE_REG_MODE = 1'b0;
defparam \LM_CK~output .OE_ASYNC_MODE = 1'b0;
defparam \LM_CK~output .OE_SYNC_MODE = 1'b0;
defparam \LM_CK~output .OE_POWERUP = 1'b0;
defparam \LM_CK~output .CFG_TRI_INPUT = 1'b0;
defparam \LM_CK~output .CFG_INPUT_EN = 1'b0;
defparam \LM_CK~output .CFG_PULL_UP = 1'b0;
defparam \LM_CK~output .CFG_SLR = 1'b0;
defparam \LM_CK~output .CFG_OPEN_DRAIN = 1'b0;
defparam \LM_CK~output .CFG_PDRCTRL = 4'b0100;
defparam \LM_CK~output .CFG_KEEP = 2'b00;
defparam \LM_CK~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \LM_CK~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \LM_CK~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \LM_CK~output .CFG_LVDS_IN_EN = 1'b0;
defparam \LM_CK~output .DPCLK_DELAY = 4'b0000;
defparam \LM_CK~output .OUT_DELAY = 1'b0;
defparam \LM_CK~output .IN_DATA_DELAY = 3'b000;
defparam \LM_CK~output .IN_REG_DELAY = 3'b000;

alta_rio \LM_D0~input (
	.padio(LM_D0),
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\LM_D0~input_o ),
	.regout());
defparam \LM_D0~input .coord_x = 16;
defparam \LM_D0~input .coord_y = 13;
defparam \LM_D0~input .coord_z = 2;
defparam \LM_D0~input .IN_ASYNC_MODE = 1'b0;
defparam \LM_D0~input .IN_SYNC_MODE = 1'b0;
defparam \LM_D0~input .IN_POWERUP = 1'b0;
defparam \LM_D0~input .OUT_REG_MODE = 1'b0;
defparam \LM_D0~input .OUT_ASYNC_MODE = 1'b0;
defparam \LM_D0~input .OUT_SYNC_MODE = 1'b0;
defparam \LM_D0~input .OUT_POWERUP = 1'b0;
defparam \LM_D0~input .OE_REG_MODE = 1'b0;
defparam \LM_D0~input .OE_ASYNC_MODE = 1'b0;
defparam \LM_D0~input .OE_SYNC_MODE = 1'b0;
defparam \LM_D0~input .OE_POWERUP = 1'b0;
defparam \LM_D0~input .CFG_TRI_INPUT = 1'b0;
defparam \LM_D0~input .CFG_INPUT_EN = 1'b1;
defparam \LM_D0~input .CFG_PULL_UP = 1'b0;
defparam \LM_D0~input .CFG_SLR = 1'b0;
defparam \LM_D0~input .CFG_OPEN_DRAIN = 1'b0;
defparam \LM_D0~input .CFG_PDRCTRL = 4'b0100;
defparam \LM_D0~input .CFG_KEEP = 2'b00;
defparam \LM_D0~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \LM_D0~input .CFG_LVDS_SEL_CUA = 2'b00;
defparam \LM_D0~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \LM_D0~input .CFG_LVDS_IN_EN = 1'b0;
defparam \LM_D0~input .DPCLK_DELAY = 4'b0000;
defparam \LM_D0~input .OUT_DELAY = 1'b0;
defparam \LM_D0~input .IN_DATA_DELAY = 3'b000;
defparam \LM_D0~input .IN_REG_DELAY = 3'b000;

alta_rio \LM_D1~input (
	.padio(LM_D1),
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\LM_D1~input_o ),
	.regout());
defparam \LM_D1~input .coord_x = 0;
defparam \LM_D1~input .coord_y = 4;
defparam \LM_D1~input .coord_z = 0;
defparam \LM_D1~input .IN_ASYNC_MODE = 1'b0;
defparam \LM_D1~input .IN_SYNC_MODE = 1'b0;
defparam \LM_D1~input .IN_POWERUP = 1'b0;
defparam \LM_D1~input .OUT_REG_MODE = 1'b0;
defparam \LM_D1~input .OUT_ASYNC_MODE = 1'b0;
defparam \LM_D1~input .OUT_SYNC_MODE = 1'b0;
defparam \LM_D1~input .OUT_POWERUP = 1'b0;
defparam \LM_D1~input .OE_REG_MODE = 1'b0;
defparam \LM_D1~input .OE_ASYNC_MODE = 1'b0;
defparam \LM_D1~input .OE_SYNC_MODE = 1'b0;
defparam \LM_D1~input .OE_POWERUP = 1'b0;
defparam \LM_D1~input .CFG_TRI_INPUT = 1'b0;
defparam \LM_D1~input .CFG_INPUT_EN = 1'b1;
defparam \LM_D1~input .CFG_PULL_UP = 1'b0;
defparam \LM_D1~input .CFG_SLR = 1'b0;
defparam \LM_D1~input .CFG_OPEN_DRAIN = 1'b0;
defparam \LM_D1~input .CFG_PDRCTRL = 4'b0100;
defparam \LM_D1~input .CFG_KEEP = 2'b00;
defparam \LM_D1~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \LM_D1~input .CFG_LVDS_SEL_CUA = 2'b00;
defparam \LM_D1~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \LM_D1~input .CFG_LVDS_IN_EN = 1'b0;
defparam \LM_D1~input .DPCLK_DELAY = 4'b0000;
defparam \LM_D1~input .OUT_DELAY = 1'b0;
defparam \LM_D1~input .IN_DATA_DELAY = 3'b000;
defparam \LM_D1~input .IN_REG_DELAY = 3'b000;

alta_rio \LM_D2~input (
	.padio(LM_D2),
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\LM_D2~input_o ),
	.regout());
defparam \LM_D2~input .coord_x = 0;
defparam \LM_D2~input .coord_y = 4;
defparam \LM_D2~input .coord_z = 3;
defparam \LM_D2~input .IN_ASYNC_MODE = 1'b0;
defparam \LM_D2~input .IN_SYNC_MODE = 1'b0;
defparam \LM_D2~input .IN_POWERUP = 1'b0;
defparam \LM_D2~input .OUT_REG_MODE = 1'b0;
defparam \LM_D2~input .OUT_ASYNC_MODE = 1'b0;
defparam \LM_D2~input .OUT_SYNC_MODE = 1'b0;
defparam \LM_D2~input .OUT_POWERUP = 1'b0;
defparam \LM_D2~input .OE_REG_MODE = 1'b0;
defparam \LM_D2~input .OE_ASYNC_MODE = 1'b0;
defparam \LM_D2~input .OE_SYNC_MODE = 1'b0;
defparam \LM_D2~input .OE_POWERUP = 1'b0;
defparam \LM_D2~input .CFG_TRI_INPUT = 1'b0;
defparam \LM_D2~input .CFG_INPUT_EN = 1'b1;
defparam \LM_D2~input .CFG_PULL_UP = 1'b0;
defparam \LM_D2~input .CFG_SLR = 1'b0;
defparam \LM_D2~input .CFG_OPEN_DRAIN = 1'b0;
defparam \LM_D2~input .CFG_PDRCTRL = 4'b0100;
defparam \LM_D2~input .CFG_KEEP = 2'b00;
defparam \LM_D2~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \LM_D2~input .CFG_LVDS_SEL_CUA = 2'b00;
defparam \LM_D2~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \LM_D2~input .CFG_LVDS_IN_EN = 1'b0;
defparam \LM_D2~input .DPCLK_DELAY = 4'b0000;
defparam \LM_D2~input .OUT_DELAY = 1'b0;
defparam \LM_D2~input .IN_DATA_DELAY = 3'b000;
defparam \LM_D2~input .IN_REG_DELAY = 3'b000;

alta_rio \LM_D3~input (
	.padio(LM_D3),
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\LM_D3~input_o ),
	.regout());
defparam \LM_D3~input .coord_x = 19;
defparam \LM_D3~input .coord_y = 0;
defparam \LM_D3~input .coord_z = 1;
defparam \LM_D3~input .IN_ASYNC_MODE = 1'b0;
defparam \LM_D3~input .IN_SYNC_MODE = 1'b0;
defparam \LM_D3~input .IN_POWERUP = 1'b0;
defparam \LM_D3~input .OUT_REG_MODE = 1'b0;
defparam \LM_D3~input .OUT_ASYNC_MODE = 1'b0;
defparam \LM_D3~input .OUT_SYNC_MODE = 1'b0;
defparam \LM_D3~input .OUT_POWERUP = 1'b0;
defparam \LM_D3~input .OE_REG_MODE = 1'b0;
defparam \LM_D3~input .OE_ASYNC_MODE = 1'b0;
defparam \LM_D3~input .OE_SYNC_MODE = 1'b0;
defparam \LM_D3~input .OE_POWERUP = 1'b0;
defparam \LM_D3~input .CFG_TRI_INPUT = 1'b0;
defparam \LM_D3~input .CFG_INPUT_EN = 1'b1;
defparam \LM_D3~input .CFG_PULL_UP = 1'b0;
defparam \LM_D3~input .CFG_SLR = 1'b0;
defparam \LM_D3~input .CFG_OPEN_DRAIN = 1'b0;
defparam \LM_D3~input .CFG_PDRCTRL = 4'b0100;
defparam \LM_D3~input .CFG_KEEP = 2'b00;
defparam \LM_D3~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \LM_D3~input .CFG_LVDS_SEL_CUA = 2'b00;
defparam \LM_D3~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \LM_D3~input .CFG_LVDS_IN_EN = 1'b0;
defparam \LM_D3~input .DPCLK_DELAY = 4'b0000;
defparam \LM_D3~input .OUT_DELAY = 1'b0;
defparam \LM_D3~input .IN_DATA_DELAY = 3'b000;
defparam \LM_D3~input .IN_REG_DELAY = 3'b000;

alta_rio \LM_D4~input (
	.padio(LM_D4),
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\LM_D4~input_o ),
	.regout());
defparam \LM_D4~input .coord_x = 22;
defparam \LM_D4~input .coord_y = 3;
defparam \LM_D4~input .coord_z = 3;
defparam \LM_D4~input .IN_ASYNC_MODE = 1'b0;
defparam \LM_D4~input .IN_SYNC_MODE = 1'b0;
defparam \LM_D4~input .IN_POWERUP = 1'b0;
defparam \LM_D4~input .OUT_REG_MODE = 1'b0;
defparam \LM_D4~input .OUT_ASYNC_MODE = 1'b0;
defparam \LM_D4~input .OUT_SYNC_MODE = 1'b0;
defparam \LM_D4~input .OUT_POWERUP = 1'b0;
defparam \LM_D4~input .OE_REG_MODE = 1'b0;
defparam \LM_D4~input .OE_ASYNC_MODE = 1'b0;
defparam \LM_D4~input .OE_SYNC_MODE = 1'b0;
defparam \LM_D4~input .OE_POWERUP = 1'b0;
defparam \LM_D4~input .CFG_TRI_INPUT = 1'b0;
defparam \LM_D4~input .CFG_INPUT_EN = 1'b1;
defparam \LM_D4~input .CFG_PULL_UP = 1'b0;
defparam \LM_D4~input .CFG_SLR = 1'b0;
defparam \LM_D4~input .CFG_OPEN_DRAIN = 1'b0;
defparam \LM_D4~input .CFG_PDRCTRL = 4'b0100;
defparam \LM_D4~input .CFG_KEEP = 2'b00;
defparam \LM_D4~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \LM_D4~input .CFG_LVDS_SEL_CUA = 2'b00;
defparam \LM_D4~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \LM_D4~input .CFG_LVDS_IN_EN = 1'b0;
defparam \LM_D4~input .DPCLK_DELAY = 4'b0000;
defparam \LM_D4~input .OUT_DELAY = 1'b0;
defparam \LM_D4~input .IN_DATA_DELAY = 3'b000;
defparam \LM_D4~input .IN_REG_DELAY = 3'b000;

alta_rio \LM_D5~input (
	.padio(LM_D5),
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\LM_D5~input_o ),
	.regout());
defparam \LM_D5~input .coord_x = 22;
defparam \LM_D5~input .coord_y = 3;
defparam \LM_D5~input .coord_z = 0;
defparam \LM_D5~input .IN_ASYNC_MODE = 1'b0;
defparam \LM_D5~input .IN_SYNC_MODE = 1'b0;
defparam \LM_D5~input .IN_POWERUP = 1'b0;
defparam \LM_D5~input .OUT_REG_MODE = 1'b0;
defparam \LM_D5~input .OUT_ASYNC_MODE = 1'b0;
defparam \LM_D5~input .OUT_SYNC_MODE = 1'b0;
defparam \LM_D5~input .OUT_POWERUP = 1'b0;
defparam \LM_D5~input .OE_REG_MODE = 1'b0;
defparam \LM_D5~input .OE_ASYNC_MODE = 1'b0;
defparam \LM_D5~input .OE_SYNC_MODE = 1'b0;
defparam \LM_D5~input .OE_POWERUP = 1'b0;
defparam \LM_D5~input .CFG_TRI_INPUT = 1'b0;
defparam \LM_D5~input .CFG_INPUT_EN = 1'b1;
defparam \LM_D5~input .CFG_PULL_UP = 1'b0;
defparam \LM_D5~input .CFG_SLR = 1'b0;
defparam \LM_D5~input .CFG_OPEN_DRAIN = 1'b0;
defparam \LM_D5~input .CFG_PDRCTRL = 4'b0100;
defparam \LM_D5~input .CFG_KEEP = 2'b00;
defparam \LM_D5~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \LM_D5~input .CFG_LVDS_SEL_CUA = 2'b00;
defparam \LM_D5~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \LM_D5~input .CFG_LVDS_IN_EN = 1'b0;
defparam \LM_D5~input .DPCLK_DELAY = 4'b0000;
defparam \LM_D5~input .OUT_DELAY = 1'b0;
defparam \LM_D5~input .IN_DATA_DELAY = 3'b000;
defparam \LM_D5~input .IN_REG_DELAY = 3'b000;

alta_rio \LM_LD~output (
	.padio(LM_LD),
	.datain(!\macro_inst|serial_lim_input_inst|load~q ),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \LM_LD~output .coord_x = 0;
defparam \LM_LD~output .coord_y = 2;
defparam \LM_LD~output .coord_z = 0;
defparam \LM_LD~output .IN_ASYNC_MODE = 1'b0;
defparam \LM_LD~output .IN_SYNC_MODE = 1'b0;
defparam \LM_LD~output .IN_POWERUP = 1'b0;
defparam \LM_LD~output .OUT_REG_MODE = 1'b0;
defparam \LM_LD~output .OUT_ASYNC_MODE = 1'b0;
defparam \LM_LD~output .OUT_SYNC_MODE = 1'b0;
defparam \LM_LD~output .OUT_POWERUP = 1'b0;
defparam \LM_LD~output .OE_REG_MODE = 1'b0;
defparam \LM_LD~output .OE_ASYNC_MODE = 1'b0;
defparam \LM_LD~output .OE_SYNC_MODE = 1'b0;
defparam \LM_LD~output .OE_POWERUP = 1'b0;
defparam \LM_LD~output .CFG_TRI_INPUT = 1'b0;
defparam \LM_LD~output .CFG_INPUT_EN = 1'b0;
defparam \LM_LD~output .CFG_PULL_UP = 1'b0;
defparam \LM_LD~output .CFG_SLR = 1'b0;
defparam \LM_LD~output .CFG_OPEN_DRAIN = 1'b0;
defparam \LM_LD~output .CFG_PDRCTRL = 4'b0100;
defparam \LM_LD~output .CFG_KEEP = 2'b00;
defparam \LM_LD~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \LM_LD~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \LM_LD~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \LM_LD~output .CFG_LVDS_IN_EN = 1'b0;
defparam \LM_LD~output .DPCLK_DELAY = 4'b0000;
defparam \LM_LD~output .OUT_DELAY = 1'b0;
defparam \LM_LD~output .IN_DATA_DELAY = 3'b000;
defparam \LM_LD~output .IN_REG_DELAY = 3'b000;

alta_rio \PIN_HSE~input (
	.padio(PIN_HSE),
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\PIN_HSE~input_o ),
	.regout());
defparam \PIN_HSE~input .coord_x = 22;
defparam \PIN_HSE~input .coord_y = 4;
defparam \PIN_HSE~input .coord_z = 1;
defparam \PIN_HSE~input .IN_ASYNC_MODE = 1'b0;
defparam \PIN_HSE~input .IN_SYNC_MODE = 1'b0;
defparam \PIN_HSE~input .IN_POWERUP = 1'b0;
defparam \PIN_HSE~input .OUT_REG_MODE = 1'b0;
defparam \PIN_HSE~input .OUT_ASYNC_MODE = 1'b0;
defparam \PIN_HSE~input .OUT_SYNC_MODE = 1'b0;
defparam \PIN_HSE~input .OUT_POWERUP = 1'b0;
defparam \PIN_HSE~input .OE_REG_MODE = 1'b0;
defparam \PIN_HSE~input .OE_ASYNC_MODE = 1'b0;
defparam \PIN_HSE~input .OE_SYNC_MODE = 1'b0;
defparam \PIN_HSE~input .OE_POWERUP = 1'b0;
defparam \PIN_HSE~input .CFG_TRI_INPUT = 1'b0;
defparam \PIN_HSE~input .CFG_PULL_UP = 1'b0;
defparam \PIN_HSE~input .CFG_SLR = 1'b0;
defparam \PIN_HSE~input .CFG_OPEN_DRAIN = 1'b0;
defparam \PIN_HSE~input .CFG_PDRCTRL = 4'b0010;
defparam \PIN_HSE~input .CFG_KEEP = 2'b00;
defparam \PIN_HSE~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \PIN_HSE~input .CFG_LVDS_SEL_CUA = 2'b00;
defparam \PIN_HSE~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \PIN_HSE~input .CFG_LVDS_IN_EN = 1'b0;
defparam \PIN_HSE~input .DPCLK_DELAY = 4'b0000;
defparam \PIN_HSE~input .OUT_DELAY = 1'b0;
defparam \PIN_HSE~input .IN_DATA_DELAY = 3'b000;
defparam \PIN_HSE~input .IN_REG_DELAY = 3'b000;

alta_rio \PIN_HSI~input (
	.padio(PIN_HSI),
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\PIN_HSI~input_o ),
	.regout());
defparam \PIN_HSI~input .coord_x = 22;
defparam \PIN_HSI~input .coord_y = 4;
defparam \PIN_HSI~input .coord_z = 0;
defparam \PIN_HSI~input .IN_ASYNC_MODE = 1'b0;
defparam \PIN_HSI~input .IN_SYNC_MODE = 1'b0;
defparam \PIN_HSI~input .IN_POWERUP = 1'b0;
defparam \PIN_HSI~input .OUT_REG_MODE = 1'b0;
defparam \PIN_HSI~input .OUT_ASYNC_MODE = 1'b0;
defparam \PIN_HSI~input .OUT_SYNC_MODE = 1'b0;
defparam \PIN_HSI~input .OUT_POWERUP = 1'b0;
defparam \PIN_HSI~input .OE_REG_MODE = 1'b0;
defparam \PIN_HSI~input .OE_ASYNC_MODE = 1'b0;
defparam \PIN_HSI~input .OE_SYNC_MODE = 1'b0;
defparam \PIN_HSI~input .OE_POWERUP = 1'b0;
defparam \PIN_HSI~input .CFG_TRI_INPUT = 1'b0;
defparam \PIN_HSI~input .CFG_PULL_UP = 1'b0;
defparam \PIN_HSI~input .CFG_SLR = 1'b0;
defparam \PIN_HSI~input .CFG_OPEN_DRAIN = 1'b0;
defparam \PIN_HSI~input .CFG_PDRCTRL = 4'b0010;
defparam \PIN_HSI~input .CFG_KEEP = 2'b00;
defparam \PIN_HSI~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \PIN_HSI~input .CFG_LVDS_SEL_CUA = 2'b00;
defparam \PIN_HSI~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \PIN_HSI~input .CFG_LVDS_IN_EN = 1'b0;
defparam \PIN_HSI~input .DPCLK_DELAY = 4'b0000;
defparam \PIN_HSI~input .OUT_DELAY = 1'b0;
defparam \PIN_HSI~input .IN_DATA_DELAY = 3'b000;
defparam \PIN_HSI~input .IN_REG_DELAY = 3'b000;

alta_rio \PIN_OSC~input (
	.padio(PIN_OSC),
	.datain(gnd),
	.oe(gnd),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(\PIN_OSC~input_o ),
	.regout());
defparam \PIN_OSC~input .coord_x = 22;
defparam \PIN_OSC~input .coord_y = 4;
defparam \PIN_OSC~input .coord_z = 2;
defparam \PIN_OSC~input .IN_ASYNC_MODE = 1'b0;
defparam \PIN_OSC~input .IN_SYNC_MODE = 1'b0;
defparam \PIN_OSC~input .IN_POWERUP = 1'b0;
defparam \PIN_OSC~input .OUT_REG_MODE = 1'b0;
defparam \PIN_OSC~input .OUT_ASYNC_MODE = 1'b0;
defparam \PIN_OSC~input .OUT_SYNC_MODE = 1'b0;
defparam \PIN_OSC~input .OUT_POWERUP = 1'b0;
defparam \PIN_OSC~input .OE_REG_MODE = 1'b0;
defparam \PIN_OSC~input .OE_ASYNC_MODE = 1'b0;
defparam \PIN_OSC~input .OE_SYNC_MODE = 1'b0;
defparam \PIN_OSC~input .OE_POWERUP = 1'b0;
defparam \PIN_OSC~input .CFG_TRI_INPUT = 1'b0;
defparam \PIN_OSC~input .CFG_PULL_UP = 1'b0;
defparam \PIN_OSC~input .CFG_SLR = 1'b0;
defparam \PIN_OSC~input .CFG_OPEN_DRAIN = 1'b0;
defparam \PIN_OSC~input .CFG_PDRCTRL = 4'b0010;
defparam \PIN_OSC~input .CFG_KEEP = 2'b00;
defparam \PIN_OSC~input .CFG_LVDS_OUT_EN = 1'b0;
defparam \PIN_OSC~input .CFG_LVDS_SEL_CUA = 2'b00;
defparam \PIN_OSC~input .CFG_LVDS_IREF = 10'b0110000000;
defparam \PIN_OSC~input .CFG_LVDS_IN_EN = 1'b0;
defparam \PIN_OSC~input .DPCLK_DELAY = 4'b0000;
defparam \PIN_OSC~input .OUT_DELAY = 1'b0;
defparam \PIN_OSC~input .IN_DATA_DELAY = 3'b000;
defparam \PIN_OSC~input .IN_REG_DELAY = 3'b000;

alta_slice PLL_ENABLE(
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.sys_ctrl_pllEnable ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\PLL_ENABLE~combout ),
	.Cout(),
	.Q());
defparam PLL_ENABLE.coord_x = 5;
defparam PLL_ENABLE.coord_y = 3;
defparam PLL_ENABLE.coord_z = 15;
defparam PLL_ENABLE.mask = 16'h00FF;
defparam PLL_ENABLE.modeMux = 1'b0;
defparam PLL_ENABLE.FeedbackMux = 1'b0;
defparam PLL_ENABLE.ShiftMux = 1'b0;
defparam PLL_ENABLE.BypassEn = 1'b0;
defparam PLL_ENABLE.CarryEnb = 1'b1;

alta_io_gclk \PLL_ENABLE~clkctrl (
	.inclk(\PLL_ENABLE~combout ),
	.outclk(\PLL_ENABLE~clkctrl_outclk ));
defparam \PLL_ENABLE~clkctrl .coord_x = 22;
defparam \PLL_ENABLE~clkctrl .coord_y = 4;
defparam \PLL_ENABLE~clkctrl .coord_z = 3;

alta_slice PLL_LOCK(
	.A(vcc),
	.B(\pll_inst|auto_generated|pll_lock_sync~q ),
	.C(vcc),
	.D(\auto_generated_inst.hbo_13_1bc039b416d3bc4a_bp ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\PLL_LOCK~combout ),
	.Cout(),
	.Q());
defparam PLL_LOCK.coord_x = 5;
defparam PLL_LOCK.coord_y = 3;
defparam PLL_LOCK.coord_z = 6;
defparam PLL_LOCK.mask = 16'hCC00;
defparam PLL_LOCK.modeMux = 1'b0;
defparam PLL_LOCK.FeedbackMux = 1'b0;
defparam PLL_LOCK.ShiftMux = 1'b0;
defparam PLL_LOCK.BypassEn = 1'b0;
defparam PLL_LOCK.CarryEnb = 1'b1;

alta_rio \SH1~output (
	.padio(SH1),
	.datain(\macro_inst|controller|serial|shi~q ),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \SH1~output .coord_x = 0;
defparam \SH1~output .coord_y = 1;
defparam \SH1~output .coord_z = 5;
defparam \SH1~output .IN_ASYNC_MODE = 1'b0;
defparam \SH1~output .IN_SYNC_MODE = 1'b0;
defparam \SH1~output .IN_POWERUP = 1'b0;
defparam \SH1~output .OUT_REG_MODE = 1'b0;
defparam \SH1~output .OUT_ASYNC_MODE = 1'b0;
defparam \SH1~output .OUT_SYNC_MODE = 1'b0;
defparam \SH1~output .OUT_POWERUP = 1'b0;
defparam \SH1~output .OE_REG_MODE = 1'b0;
defparam \SH1~output .OE_ASYNC_MODE = 1'b0;
defparam \SH1~output .OE_SYNC_MODE = 1'b0;
defparam \SH1~output .OE_POWERUP = 1'b0;
defparam \SH1~output .CFG_TRI_INPUT = 1'b0;
defparam \SH1~output .CFG_INPUT_EN = 1'b0;
defparam \SH1~output .CFG_PULL_UP = 1'b0;
defparam \SH1~output .CFG_SLR = 1'b0;
defparam \SH1~output .CFG_OPEN_DRAIN = 1'b0;
defparam \SH1~output .CFG_PDRCTRL = 4'b0100;
defparam \SH1~output .CFG_KEEP = 2'b00;
defparam \SH1~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \SH1~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \SH1~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \SH1~output .CFG_LVDS_IN_EN = 1'b0;
defparam \SH1~output .DPCLK_DELAY = 4'b0000;
defparam \SH1~output .OUT_DELAY = 1'b0;
defparam \SH1~output .IN_DATA_DELAY = 3'b000;
defparam \SH1~output .IN_REG_DELAY = 3'b000;

alta_rio \SH2~output (
	.padio(SH2),
	.datain(\macro_inst|controller|serial|shi~q ),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \SH2~output .coord_x = 0;
defparam \SH2~output .coord_y = 1;
defparam \SH2~output .coord_z = 0;
defparam \SH2~output .IN_ASYNC_MODE = 1'b0;
defparam \SH2~output .IN_SYNC_MODE = 1'b0;
defparam \SH2~output .IN_POWERUP = 1'b0;
defparam \SH2~output .OUT_REG_MODE = 1'b0;
defparam \SH2~output .OUT_ASYNC_MODE = 1'b0;
defparam \SH2~output .OUT_SYNC_MODE = 1'b0;
defparam \SH2~output .OUT_POWERUP = 1'b0;
defparam \SH2~output .OE_REG_MODE = 1'b0;
defparam \SH2~output .OE_ASYNC_MODE = 1'b0;
defparam \SH2~output .OE_SYNC_MODE = 1'b0;
defparam \SH2~output .OE_POWERUP = 1'b0;
defparam \SH2~output .CFG_TRI_INPUT = 1'b0;
defparam \SH2~output .CFG_INPUT_EN = 1'b0;
defparam \SH2~output .CFG_PULL_UP = 1'b0;
defparam \SH2~output .CFG_SLR = 1'b0;
defparam \SH2~output .CFG_OPEN_DRAIN = 1'b0;
defparam \SH2~output .CFG_PDRCTRL = 4'b0100;
defparam \SH2~output .CFG_KEEP = 2'b00;
defparam \SH2~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \SH2~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \SH2~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \SH2~output .CFG_LVDS_IN_EN = 1'b0;
defparam \SH2~output .DPCLK_DELAY = 4'b0000;
defparam \SH2~output .OUT_DELAY = 1'b0;
defparam \SH2~output .IN_DATA_DELAY = 3'b000;
defparam \SH2~output .IN_REG_DELAY = 3'b000;

alta_rio \SH3~output (
	.padio(SH3),
	.datain(\macro_inst|controller|serial|shi~q ),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \SH3~output .coord_x = 0;
defparam \SH3~output .coord_y = 2;
defparam \SH3~output .coord_z = 3;
defparam \SH3~output .IN_ASYNC_MODE = 1'b0;
defparam \SH3~output .IN_SYNC_MODE = 1'b0;
defparam \SH3~output .IN_POWERUP = 1'b0;
defparam \SH3~output .OUT_REG_MODE = 1'b0;
defparam \SH3~output .OUT_ASYNC_MODE = 1'b0;
defparam \SH3~output .OUT_SYNC_MODE = 1'b0;
defparam \SH3~output .OUT_POWERUP = 1'b0;
defparam \SH3~output .OE_REG_MODE = 1'b0;
defparam \SH3~output .OE_ASYNC_MODE = 1'b0;
defparam \SH3~output .OE_SYNC_MODE = 1'b0;
defparam \SH3~output .OE_POWERUP = 1'b0;
defparam \SH3~output .CFG_TRI_INPUT = 1'b0;
defparam \SH3~output .CFG_INPUT_EN = 1'b0;
defparam \SH3~output .CFG_PULL_UP = 1'b0;
defparam \SH3~output .CFG_SLR = 1'b0;
defparam \SH3~output .CFG_OPEN_DRAIN = 1'b0;
defparam \SH3~output .CFG_PDRCTRL = 4'b0100;
defparam \SH3~output .CFG_KEEP = 2'b00;
defparam \SH3~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \SH3~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \SH3~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \SH3~output .CFG_LVDS_IN_EN = 1'b0;
defparam \SH3~output .DPCLK_DELAY = 4'b0000;
defparam \SH3~output .OUT_DELAY = 1'b0;
defparam \SH3~output .IN_DATA_DELAY = 3'b000;
defparam \SH3~output .IN_REG_DELAY = 3'b000;

alta_rio \SH4~output (
	.padio(SH4),
	.datain(\macro_inst|controller|serial|shi~q ),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \SH4~output .coord_x = 18;
defparam \SH4~output .coord_y = 13;
defparam \SH4~output .coord_z = 3;
defparam \SH4~output .IN_ASYNC_MODE = 1'b0;
defparam \SH4~output .IN_SYNC_MODE = 1'b0;
defparam \SH4~output .IN_POWERUP = 1'b0;
defparam \SH4~output .OUT_REG_MODE = 1'b0;
defparam \SH4~output .OUT_ASYNC_MODE = 1'b0;
defparam \SH4~output .OUT_SYNC_MODE = 1'b0;
defparam \SH4~output .OUT_POWERUP = 1'b0;
defparam \SH4~output .OE_REG_MODE = 1'b0;
defparam \SH4~output .OE_ASYNC_MODE = 1'b0;
defparam \SH4~output .OE_SYNC_MODE = 1'b0;
defparam \SH4~output .OE_POWERUP = 1'b0;
defparam \SH4~output .CFG_TRI_INPUT = 1'b0;
defparam \SH4~output .CFG_INPUT_EN = 1'b0;
defparam \SH4~output .CFG_PULL_UP = 1'b0;
defparam \SH4~output .CFG_SLR = 1'b0;
defparam \SH4~output .CFG_OPEN_DRAIN = 1'b0;
defparam \SH4~output .CFG_PDRCTRL = 4'b0100;
defparam \SH4~output .CFG_KEEP = 2'b00;
defparam \SH4~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \SH4~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \SH4~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \SH4~output .CFG_LVDS_IN_EN = 1'b0;
defparam \SH4~output .DPCLK_DELAY = 4'b0000;
defparam \SH4~output .OUT_DELAY = 1'b0;
defparam \SH4~output .IN_DATA_DELAY = 3'b000;
defparam \SH4~output .IN_REG_DELAY = 3'b000;

alta_rio \SH5~output (
	.padio(SH5),
	.datain(\macro_inst|controller|serial|shi~q ),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \SH5~output .coord_x = 19;
defparam \SH5~output .coord_y = 13;
defparam \SH5~output .coord_z = 2;
defparam \SH5~output .IN_ASYNC_MODE = 1'b0;
defparam \SH5~output .IN_SYNC_MODE = 1'b0;
defparam \SH5~output .IN_POWERUP = 1'b0;
defparam \SH5~output .OUT_REG_MODE = 1'b0;
defparam \SH5~output .OUT_ASYNC_MODE = 1'b0;
defparam \SH5~output .OUT_SYNC_MODE = 1'b0;
defparam \SH5~output .OUT_POWERUP = 1'b0;
defparam \SH5~output .OE_REG_MODE = 1'b0;
defparam \SH5~output .OE_ASYNC_MODE = 1'b0;
defparam \SH5~output .OE_SYNC_MODE = 1'b0;
defparam \SH5~output .OE_POWERUP = 1'b0;
defparam \SH5~output .CFG_TRI_INPUT = 1'b0;
defparam \SH5~output .CFG_INPUT_EN = 1'b0;
defparam \SH5~output .CFG_PULL_UP = 1'b0;
defparam \SH5~output .CFG_SLR = 1'b0;
defparam \SH5~output .CFG_OPEN_DRAIN = 1'b0;
defparam \SH5~output .CFG_PDRCTRL = 4'b0100;
defparam \SH5~output .CFG_KEEP = 2'b00;
defparam \SH5~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \SH5~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \SH5~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \SH5~output .CFG_LVDS_IN_EN = 1'b0;
defparam \SH5~output .DPCLK_DELAY = 4'b0000;
defparam \SH5~output .OUT_DELAY = 1'b0;
defparam \SH5~output .IN_DATA_DELAY = 3'b000;
defparam \SH5~output .IN_REG_DELAY = 3'b000;

alta_rio \SH6~output (
	.padio(SH6),
	.datain(\macro_inst|controller|serial|shi~q ),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \SH6~output .coord_x = 20;
defparam \SH6~output .coord_y = 13;
defparam \SH6~output .coord_z = 2;
defparam \SH6~output .IN_ASYNC_MODE = 1'b0;
defparam \SH6~output .IN_SYNC_MODE = 1'b0;
defparam \SH6~output .IN_POWERUP = 1'b0;
defparam \SH6~output .OUT_REG_MODE = 1'b0;
defparam \SH6~output .OUT_ASYNC_MODE = 1'b0;
defparam \SH6~output .OUT_SYNC_MODE = 1'b0;
defparam \SH6~output .OUT_POWERUP = 1'b0;
defparam \SH6~output .OE_REG_MODE = 1'b0;
defparam \SH6~output .OE_ASYNC_MODE = 1'b0;
defparam \SH6~output .OE_SYNC_MODE = 1'b0;
defparam \SH6~output .OE_POWERUP = 1'b0;
defparam \SH6~output .CFG_TRI_INPUT = 1'b0;
defparam \SH6~output .CFG_INPUT_EN = 1'b0;
defparam \SH6~output .CFG_PULL_UP = 1'b0;
defparam \SH6~output .CFG_SLR = 1'b0;
defparam \SH6~output .CFG_OPEN_DRAIN = 1'b0;
defparam \SH6~output .CFG_PDRCTRL = 4'b0100;
defparam \SH6~output .CFG_KEEP = 2'b00;
defparam \SH6~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \SH6~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \SH6~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \SH6~output .CFG_LVDS_IN_EN = 1'b0;
defparam \SH6~output .DPCLK_DELAY = 4'b0000;
defparam \SH6~output .OUT_DELAY = 1'b0;
defparam \SH6~output .IN_DATA_DELAY = 3'b000;
defparam \SH6~output .IN_REG_DELAY = 3'b000;

alta_rio \ST1~output (
	.padio(ST1),
	.datain(\macro_inst|controller|serial|sto~q ),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \ST1~output .coord_x = 0;
defparam \ST1~output .coord_y = 2;
defparam \ST1~output .coord_z = 2;
defparam \ST1~output .IN_ASYNC_MODE = 1'b0;
defparam \ST1~output .IN_SYNC_MODE = 1'b0;
defparam \ST1~output .IN_POWERUP = 1'b0;
defparam \ST1~output .OUT_REG_MODE = 1'b0;
defparam \ST1~output .OUT_ASYNC_MODE = 1'b0;
defparam \ST1~output .OUT_SYNC_MODE = 1'b0;
defparam \ST1~output .OUT_POWERUP = 1'b0;
defparam \ST1~output .OE_REG_MODE = 1'b0;
defparam \ST1~output .OE_ASYNC_MODE = 1'b0;
defparam \ST1~output .OE_SYNC_MODE = 1'b0;
defparam \ST1~output .OE_POWERUP = 1'b0;
defparam \ST1~output .CFG_TRI_INPUT = 1'b0;
defparam \ST1~output .CFG_INPUT_EN = 1'b0;
defparam \ST1~output .CFG_PULL_UP = 1'b0;
defparam \ST1~output .CFG_SLR = 1'b0;
defparam \ST1~output .CFG_OPEN_DRAIN = 1'b0;
defparam \ST1~output .CFG_PDRCTRL = 4'b0100;
defparam \ST1~output .CFG_KEEP = 2'b00;
defparam \ST1~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \ST1~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \ST1~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \ST1~output .CFG_LVDS_IN_EN = 1'b0;
defparam \ST1~output .DPCLK_DELAY = 4'b0000;
defparam \ST1~output .OUT_DELAY = 1'b0;
defparam \ST1~output .IN_DATA_DELAY = 3'b000;
defparam \ST1~output .IN_REG_DELAY = 3'b000;

alta_rio \ST2~output (
	.padio(ST2),
	.datain(\macro_inst|controller|serial|sto~q ),
	.oe(vcc),
	.outclk(gnd),
	.outclkena(vcc),
	.inclk(gnd),
	.inclkena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.combout(),
	.regout());
defparam \ST2~output .coord_x = 20;
defparam \ST2~output .coord_y = 13;
defparam \ST2~output .coord_z = 1;
defparam \ST2~output .IN_ASYNC_MODE = 1'b0;
defparam \ST2~output .IN_SYNC_MODE = 1'b0;
defparam \ST2~output .IN_POWERUP = 1'b0;
defparam \ST2~output .OUT_REG_MODE = 1'b0;
defparam \ST2~output .OUT_ASYNC_MODE = 1'b0;
defparam \ST2~output .OUT_SYNC_MODE = 1'b0;
defparam \ST2~output .OUT_POWERUP = 1'b0;
defparam \ST2~output .OE_REG_MODE = 1'b0;
defparam \ST2~output .OE_ASYNC_MODE = 1'b0;
defparam \ST2~output .OE_SYNC_MODE = 1'b0;
defparam \ST2~output .OE_POWERUP = 1'b0;
defparam \ST2~output .CFG_TRI_INPUT = 1'b0;
defparam \ST2~output .CFG_INPUT_EN = 1'b0;
defparam \ST2~output .CFG_PULL_UP = 1'b0;
defparam \ST2~output .CFG_SLR = 1'b0;
defparam \ST2~output .CFG_OPEN_DRAIN = 1'b0;
defparam \ST2~output .CFG_PDRCTRL = 4'b0100;
defparam \ST2~output .CFG_KEEP = 2'b00;
defparam \ST2~output .CFG_LVDS_OUT_EN = 1'b0;
defparam \ST2~output .CFG_LVDS_SEL_CUA = 2'b00;
defparam \ST2~output .CFG_LVDS_IREF = 10'b0110000000;
defparam \ST2~output .CFG_LVDS_IN_EN = 1'b0;
defparam \ST2~output .DPCLK_DELAY = 4'b0000;
defparam \ST2~output .OUT_DELAY = 1'b0;
defparam \ST2~output .IN_DATA_DELAY = 3'b000;
defparam \ST2~output .IN_REG_DELAY = 3'b000;

alta_asyncctrl asyncreset_ctrl_X43_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ));
defparam asyncreset_ctrl_X43_Y2_N0.coord_x = 7;
defparam asyncreset_ctrl_X43_Y2_N0.coord_y = 2;
defparam asyncreset_ctrl_X43_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X43_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X46_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ));
defparam asyncreset_ctrl_X46_Y2_N0.coord_x = 4;
defparam asyncreset_ctrl_X46_Y2_N0.coord_y = 3;
defparam asyncreset_ctrl_X46_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X46_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X46_Y3_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y3_SIG ));
defparam asyncreset_ctrl_X46_Y3_N0.coord_x = 5;
defparam asyncreset_ctrl_X46_Y3_N0.coord_y = 4;
defparam asyncreset_ctrl_X46_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X46_Y3_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X47_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X47_Y2_SIG ));
defparam asyncreset_ctrl_X47_Y2_N0.coord_x = 4;
defparam asyncreset_ctrl_X47_Y2_N0.coord_y = 2;
defparam asyncreset_ctrl_X47_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X47_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X47_Y3_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X47_Y3_SIG ));
defparam asyncreset_ctrl_X47_Y3_N0.coord_x = 4;
defparam asyncreset_ctrl_X47_Y3_N0.coord_y = 4;
defparam asyncreset_ctrl_X47_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X47_Y3_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X48_Y1_N0(
	.Din(\PLL_ENABLE~clkctrl_outclk ),
	.Dout(\PLL_ENABLE~clkctrl_outclk__AsyncReset_X48_Y1_SIG ));
defparam asyncreset_ctrl_X48_Y1_N0.coord_x = 5;
defparam asyncreset_ctrl_X48_Y1_N0.coord_y = 3;
defparam asyncreset_ctrl_X48_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X48_Y1_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X48_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y2_SIG ));
defparam asyncreset_ctrl_X48_Y2_N0.coord_x = 3;
defparam asyncreset_ctrl_X48_Y2_N0.coord_y = 1;
defparam asyncreset_ctrl_X48_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X48_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X48_Y3_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y3_SIG ));
defparam asyncreset_ctrl_X48_Y3_N0.coord_x = 3;
defparam asyncreset_ctrl_X48_Y3_N0.coord_y = 2;
defparam asyncreset_ctrl_X48_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X48_Y3_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X49_Y1_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y1_SIG ));
defparam asyncreset_ctrl_X49_Y1_N0.coord_x = 6;
defparam asyncreset_ctrl_X49_Y1_N0.coord_y = 1;
defparam asyncreset_ctrl_X49_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X49_Y1_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X49_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y2_SIG ));
defparam asyncreset_ctrl_X49_Y2_N0.coord_x = 9;
defparam asyncreset_ctrl_X49_Y2_N0.coord_y = 3;
defparam asyncreset_ctrl_X49_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X49_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X49_Y2_N1(
	.Din(),
	.Dout(AsyncReset_X49_Y2_GND));
defparam asyncreset_ctrl_X49_Y2_N1.coord_x = 9;
defparam asyncreset_ctrl_X49_Y2_N1.coord_y = 3;
defparam asyncreset_ctrl_X49_Y2_N1.coord_z = 1;
defparam asyncreset_ctrl_X49_Y2_N1.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X49_Y3_N0(
	.Din(),
	.Dout(AsyncReset_X49_Y3_GND));
defparam asyncreset_ctrl_X49_Y3_N0.coord_x = 6;
defparam asyncreset_ctrl_X49_Y3_N0.coord_y = 4;
defparam asyncreset_ctrl_X49_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X49_Y3_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X49_Y4_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y4_SIG ));
defparam asyncreset_ctrl_X49_Y4_N0.coord_x = 3;
defparam asyncreset_ctrl_X49_Y4_N0.coord_y = 4;
defparam asyncreset_ctrl_X49_Y4_N0.coord_z = 0;
defparam asyncreset_ctrl_X49_Y4_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X50_Y1_N1(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y1_SIG ));
defparam asyncreset_ctrl_X50_Y1_N1.coord_x = 7;
defparam asyncreset_ctrl_X50_Y1_N1.coord_y = 1;
defparam asyncreset_ctrl_X50_Y1_N1.coord_z = 1;
defparam asyncreset_ctrl_X50_Y1_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X50_Y2_N1(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y2_SIG ));
defparam asyncreset_ctrl_X50_Y2_N1.coord_x = 9;
defparam asyncreset_ctrl_X50_Y2_N1.coord_y = 2;
defparam asyncreset_ctrl_X50_Y2_N1.coord_z = 1;
defparam asyncreset_ctrl_X50_Y2_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X50_Y3_N0(
	.Din(),
	.Dout(AsyncReset_X50_Y3_GND));
defparam asyncreset_ctrl_X50_Y3_N0.coord_x = 8;
defparam asyncreset_ctrl_X50_Y3_N0.coord_y = 4;
defparam asyncreset_ctrl_X50_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X50_Y3_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X50_Y4_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y4_SIG ));
defparam asyncreset_ctrl_X50_Y4_N0.coord_x = 9;
defparam asyncreset_ctrl_X50_Y4_N0.coord_y = 1;
defparam asyncreset_ctrl_X50_Y4_N0.coord_z = 0;
defparam asyncreset_ctrl_X50_Y4_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X51_Y1_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y1_SIG ));
defparam asyncreset_ctrl_X51_Y1_N0.coord_x = 8;
defparam asyncreset_ctrl_X51_Y1_N0.coord_y = 1;
defparam asyncreset_ctrl_X51_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X51_Y1_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X51_Y2_N1(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y2_SIG ));
defparam asyncreset_ctrl_X51_Y2_N1.coord_x = 8;
defparam asyncreset_ctrl_X51_Y2_N1.coord_y = 2;
defparam asyncreset_ctrl_X51_Y2_N1.coord_z = 1;
defparam asyncreset_ctrl_X51_Y2_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X51_Y3_N0(
	.Din(),
	.Dout(AsyncReset_X51_Y3_GND));
defparam asyncreset_ctrl_X51_Y3_N0.coord_x = 9;
defparam asyncreset_ctrl_X51_Y3_N0.coord_y = 4;
defparam asyncreset_ctrl_X51_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X51_Y3_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X51_Y3_N1(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y3_SIG ));
defparam asyncreset_ctrl_X51_Y3_N1.coord_x = 9;
defparam asyncreset_ctrl_X51_Y3_N1.coord_y = 4;
defparam asyncreset_ctrl_X51_Y3_N1.coord_z = 1;
defparam asyncreset_ctrl_X51_Y3_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X51_Y4_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ));
defparam asyncreset_ctrl_X51_Y4_N0.coord_x = 15;
defparam asyncreset_ctrl_X51_Y4_N0.coord_y = 2;
defparam asyncreset_ctrl_X51_Y4_N0.coord_z = 0;
defparam asyncreset_ctrl_X51_Y4_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X52_Y1_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ));
defparam asyncreset_ctrl_X52_Y1_N0.coord_x = 11;
defparam asyncreset_ctrl_X52_Y1_N0.coord_y = 1;
defparam asyncreset_ctrl_X52_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X52_Y1_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X52_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ));
defparam asyncreset_ctrl_X52_Y2_N0.coord_x = 16;
defparam asyncreset_ctrl_X52_Y2_N0.coord_y = 5;
defparam asyncreset_ctrl_X52_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X52_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X52_Y3_N0(
	.Din(),
	.Dout(AsyncReset_X52_Y3_GND));
defparam asyncreset_ctrl_X52_Y3_N0.coord_x = 8;
defparam asyncreset_ctrl_X52_Y3_N0.coord_y = 3;
defparam asyncreset_ctrl_X52_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X52_Y3_N0.AsyncCtrlMux = 2'b00;

alta_asyncctrl asyncreset_ctrl_X52_Y4_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ));
defparam asyncreset_ctrl_X52_Y4_N0.coord_x = 16;
defparam asyncreset_ctrl_X52_Y4_N0.coord_y = 2;
defparam asyncreset_ctrl_X52_Y4_N0.coord_z = 0;
defparam asyncreset_ctrl_X52_Y4_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X53_Y1_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ));
defparam asyncreset_ctrl_X53_Y1_N0.coord_x = 16;
defparam asyncreset_ctrl_X53_Y1_N0.coord_y = 1;
defparam asyncreset_ctrl_X53_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X53_Y1_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X53_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ));
defparam asyncreset_ctrl_X53_Y2_N0.coord_x = 19;
defparam asyncreset_ctrl_X53_Y2_N0.coord_y = 5;
defparam asyncreset_ctrl_X53_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X53_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X53_Y3_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ));
defparam asyncreset_ctrl_X53_Y3_N0.coord_x = 7;
defparam asyncreset_ctrl_X53_Y3_N0.coord_y = 4;
defparam asyncreset_ctrl_X53_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X53_Y3_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X53_Y4_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ));
defparam asyncreset_ctrl_X53_Y4_N0.coord_x = 15;
defparam asyncreset_ctrl_X53_Y4_N0.coord_y = 4;
defparam asyncreset_ctrl_X53_Y4_N0.coord_z = 0;
defparam asyncreset_ctrl_X53_Y4_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X54_Y1_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ));
defparam asyncreset_ctrl_X54_Y1_N0.coord_x = 20;
defparam asyncreset_ctrl_X54_Y1_N0.coord_y = 2;
defparam asyncreset_ctrl_X54_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X54_Y1_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X54_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y2_SIG ));
defparam asyncreset_ctrl_X54_Y2_N0.coord_x = 14;
defparam asyncreset_ctrl_X54_Y2_N0.coord_y = 5;
defparam asyncreset_ctrl_X54_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X54_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X54_Y3_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ));
defparam asyncreset_ctrl_X54_Y3_N0.coord_x = 14;
defparam asyncreset_ctrl_X54_Y3_N0.coord_y = 12;
defparam asyncreset_ctrl_X54_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X54_Y3_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X54_Y4_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ));
defparam asyncreset_ctrl_X54_Y4_N0.coord_x = 11;
defparam asyncreset_ctrl_X54_Y4_N0.coord_y = 2;
defparam asyncreset_ctrl_X54_Y4_N0.coord_z = 0;
defparam asyncreset_ctrl_X54_Y4_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X56_Y10_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ));
defparam asyncreset_ctrl_X56_Y10_N0.coord_x = 11;
defparam asyncreset_ctrl_X56_Y10_N0.coord_y = 3;
defparam asyncreset_ctrl_X56_Y10_N0.coord_z = 0;
defparam asyncreset_ctrl_X56_Y10_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X56_Y11_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ));
defparam asyncreset_ctrl_X56_Y11_N0.coord_x = 19;
defparam asyncreset_ctrl_X56_Y11_N0.coord_y = 10;
defparam asyncreset_ctrl_X56_Y11_N0.coord_z = 0;
defparam asyncreset_ctrl_X56_Y11_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X56_Y12_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ));
defparam asyncreset_ctrl_X56_Y12_N0.coord_x = 20;
defparam asyncreset_ctrl_X56_Y12_N0.coord_y = 8;
defparam asyncreset_ctrl_X56_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X56_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X56_Y1_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ));
defparam asyncreset_ctrl_X56_Y1_N0.coord_x = 10;
defparam asyncreset_ctrl_X56_Y1_N0.coord_y = 2;
defparam asyncreset_ctrl_X56_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X56_Y1_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X56_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y2_SIG ));
defparam asyncreset_ctrl_X56_Y2_N0.coord_x = 16;
defparam asyncreset_ctrl_X56_Y2_N0.coord_y = 11;
defparam asyncreset_ctrl_X56_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X56_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X56_Y3_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ));
defparam asyncreset_ctrl_X56_Y3_N0.coord_x = 12;
defparam asyncreset_ctrl_X56_Y3_N0.coord_y = 4;
defparam asyncreset_ctrl_X56_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X56_Y3_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X56_Y4_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ));
defparam asyncreset_ctrl_X56_Y4_N0.coord_x = 17;
defparam asyncreset_ctrl_X56_Y4_N0.coord_y = 4;
defparam asyncreset_ctrl_X56_Y4_N0.coord_z = 0;
defparam asyncreset_ctrl_X56_Y4_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X56_Y5_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ));
defparam asyncreset_ctrl_X56_Y5_N0.coord_x = 10;
defparam asyncreset_ctrl_X56_Y5_N0.coord_y = 4;
defparam asyncreset_ctrl_X56_Y5_N0.coord_z = 0;
defparam asyncreset_ctrl_X56_Y5_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X56_Y6_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ));
defparam asyncreset_ctrl_X56_Y6_N0.coord_x = 17;
defparam asyncreset_ctrl_X56_Y6_N0.coord_y = 2;
defparam asyncreset_ctrl_X56_Y6_N0.coord_z = 0;
defparam asyncreset_ctrl_X56_Y6_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X56_Y7_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ));
defparam asyncreset_ctrl_X56_Y7_N0.coord_x = 14;
defparam asyncreset_ctrl_X56_Y7_N0.coord_y = 2;
defparam asyncreset_ctrl_X56_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X56_Y7_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X56_Y8_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ));
defparam asyncreset_ctrl_X56_Y8_N0.coord_x = 19;
defparam asyncreset_ctrl_X56_Y8_N0.coord_y = 1;
defparam asyncreset_ctrl_X56_Y8_N0.coord_z = 0;
defparam asyncreset_ctrl_X56_Y8_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X56_Y9_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y9_SIG ));
defparam asyncreset_ctrl_X56_Y9_N0.coord_x = 17;
defparam asyncreset_ctrl_X56_Y9_N0.coord_y = 9;
defparam asyncreset_ctrl_X56_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X56_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X57_Y10_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ));
defparam asyncreset_ctrl_X57_Y10_N0.coord_x = 12;
defparam asyncreset_ctrl_X57_Y10_N0.coord_y = 3;
defparam asyncreset_ctrl_X57_Y10_N0.coord_z = 0;
defparam asyncreset_ctrl_X57_Y10_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X57_Y11_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ));
defparam asyncreset_ctrl_X57_Y11_N0.coord_x = 20;
defparam asyncreset_ctrl_X57_Y11_N0.coord_y = 10;
defparam asyncreset_ctrl_X57_Y11_N0.coord_z = 0;
defparam asyncreset_ctrl_X57_Y11_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X57_Y12_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y12_SIG ));
defparam asyncreset_ctrl_X57_Y12_N0.coord_x = 18;
defparam asyncreset_ctrl_X57_Y12_N0.coord_y = 8;
defparam asyncreset_ctrl_X57_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X57_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X57_Y1_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y1_SIG ));
defparam asyncreset_ctrl_X57_Y1_N0.coord_x = 12;
defparam asyncreset_ctrl_X57_Y1_N0.coord_y = 2;
defparam asyncreset_ctrl_X57_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X57_Y1_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X57_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ));
defparam asyncreset_ctrl_X57_Y2_N0.coord_x = 18;
defparam asyncreset_ctrl_X57_Y2_N0.coord_y = 12;
defparam asyncreset_ctrl_X57_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X57_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X57_Y3_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y3_SIG ));
defparam asyncreset_ctrl_X57_Y3_N0.coord_x = 14;
defparam asyncreset_ctrl_X57_Y3_N0.coord_y = 11;
defparam asyncreset_ctrl_X57_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X57_Y3_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X57_Y4_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ));
defparam asyncreset_ctrl_X57_Y4_N0.coord_x = 16;
defparam asyncreset_ctrl_X57_Y4_N0.coord_y = 4;
defparam asyncreset_ctrl_X57_Y4_N0.coord_z = 0;
defparam asyncreset_ctrl_X57_Y4_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X57_Y5_N1(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y5_SIG ));
defparam asyncreset_ctrl_X57_Y5_N1.coord_x = 14;
defparam asyncreset_ctrl_X57_Y5_N1.coord_y = 7;
defparam asyncreset_ctrl_X57_Y5_N1.coord_z = 1;
defparam asyncreset_ctrl_X57_Y5_N1.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X57_Y6_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y6_SIG ));
defparam asyncreset_ctrl_X57_Y6_N0.coord_x = 14;
defparam asyncreset_ctrl_X57_Y6_N0.coord_y = 10;
defparam asyncreset_ctrl_X57_Y6_N0.coord_z = 0;
defparam asyncreset_ctrl_X57_Y6_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X57_Y7_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ));
defparam asyncreset_ctrl_X57_Y7_N0.coord_x = 15;
defparam asyncreset_ctrl_X57_Y7_N0.coord_y = 3;
defparam asyncreset_ctrl_X57_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X57_Y7_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X57_Y8_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y8_SIG ));
defparam asyncreset_ctrl_X57_Y8_N0.coord_x = 18;
defparam asyncreset_ctrl_X57_Y8_N0.coord_y = 3;
defparam asyncreset_ctrl_X57_Y8_N0.coord_z = 0;
defparam asyncreset_ctrl_X57_Y8_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X57_Y9_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ));
defparam asyncreset_ctrl_X57_Y9_N0.coord_x = 16;
defparam asyncreset_ctrl_X57_Y9_N0.coord_y = 9;
defparam asyncreset_ctrl_X57_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X57_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X58_Y10_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y10_SIG ));
defparam asyncreset_ctrl_X58_Y10_N0.coord_x = 17;
defparam asyncreset_ctrl_X58_Y10_N0.coord_y = 7;
defparam asyncreset_ctrl_X58_Y10_N0.coord_z = 0;
defparam asyncreset_ctrl_X58_Y10_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X58_Y11_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ));
defparam asyncreset_ctrl_X58_Y11_N0.coord_x = 19;
defparam asyncreset_ctrl_X58_Y11_N0.coord_y = 12;
defparam asyncreset_ctrl_X58_Y11_N0.coord_z = 0;
defparam asyncreset_ctrl_X58_Y11_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X58_Y12_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y12_SIG ));
defparam asyncreset_ctrl_X58_Y12_N0.coord_x = 20;
defparam asyncreset_ctrl_X58_Y12_N0.coord_y = 3;
defparam asyncreset_ctrl_X58_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X58_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X58_Y1_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ));
defparam asyncreset_ctrl_X58_Y1_N0.coord_x = 10;
defparam asyncreset_ctrl_X58_Y1_N0.coord_y = 1;
defparam asyncreset_ctrl_X58_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X58_Y1_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X58_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ));
defparam asyncreset_ctrl_X58_Y2_N0.coord_x = 16;
defparam asyncreset_ctrl_X58_Y2_N0.coord_y = 10;
defparam asyncreset_ctrl_X58_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X58_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X58_Y3_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y3_SIG ));
defparam asyncreset_ctrl_X58_Y3_N0.coord_x = 15;
defparam asyncreset_ctrl_X58_Y3_N0.coord_y = 11;
defparam asyncreset_ctrl_X58_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X58_Y3_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X58_Y4_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y4_SIG ));
defparam asyncreset_ctrl_X58_Y4_N0.coord_x = 16;
defparam asyncreset_ctrl_X58_Y4_N0.coord_y = 8;
defparam asyncreset_ctrl_X58_Y4_N0.coord_z = 0;
defparam asyncreset_ctrl_X58_Y4_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X58_Y5_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y5_SIG ));
defparam asyncreset_ctrl_X58_Y5_N0.coord_x = 16;
defparam asyncreset_ctrl_X58_Y5_N0.coord_y = 12;
defparam asyncreset_ctrl_X58_Y5_N0.coord_z = 0;
defparam asyncreset_ctrl_X58_Y5_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X58_Y6_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ));
defparam asyncreset_ctrl_X58_Y6_N0.coord_x = 14;
defparam asyncreset_ctrl_X58_Y6_N0.coord_y = 9;
defparam asyncreset_ctrl_X58_Y6_N0.coord_z = 0;
defparam asyncreset_ctrl_X58_Y6_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X58_Y7_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y7_SIG ));
defparam asyncreset_ctrl_X58_Y7_N0.coord_x = 14;
defparam asyncreset_ctrl_X58_Y7_N0.coord_y = 4;
defparam asyncreset_ctrl_X58_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X58_Y7_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X58_Y8_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y8_SIG ));
defparam asyncreset_ctrl_X58_Y8_N0.coord_x = 17;
defparam asyncreset_ctrl_X58_Y8_N0.coord_y = 5;
defparam asyncreset_ctrl_X58_Y8_N0.coord_z = 0;
defparam asyncreset_ctrl_X58_Y8_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X58_Y9_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ));
defparam asyncreset_ctrl_X58_Y9_N0.coord_x = 18;
defparam asyncreset_ctrl_X58_Y9_N0.coord_y = 9;
defparam asyncreset_ctrl_X58_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X58_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X59_Y10_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ));
defparam asyncreset_ctrl_X59_Y10_N0.coord_x = 18;
defparam asyncreset_ctrl_X59_Y10_N0.coord_y = 6;
defparam asyncreset_ctrl_X59_Y10_N0.coord_z = 0;
defparam asyncreset_ctrl_X59_Y10_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X59_Y11_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y11_SIG ));
defparam asyncreset_ctrl_X59_Y11_N0.coord_x = 19;
defparam asyncreset_ctrl_X59_Y11_N0.coord_y = 3;
defparam asyncreset_ctrl_X59_Y11_N0.coord_z = 0;
defparam asyncreset_ctrl_X59_Y11_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X59_Y12_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ));
defparam asyncreset_ctrl_X59_Y12_N0.coord_x = 20;
defparam asyncreset_ctrl_X59_Y12_N0.coord_y = 5;
defparam asyncreset_ctrl_X59_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X59_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X59_Y1_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ));
defparam asyncreset_ctrl_X59_Y1_N0.coord_x = 16;
defparam asyncreset_ctrl_X59_Y1_N0.coord_y = 3;
defparam asyncreset_ctrl_X59_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X59_Y1_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X59_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ));
defparam asyncreset_ctrl_X59_Y2_N0.coord_x = 10;
defparam asyncreset_ctrl_X59_Y2_N0.coord_y = 3;
defparam asyncreset_ctrl_X59_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X59_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X59_Y3_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y3_SIG ));
defparam asyncreset_ctrl_X59_Y3_N0.coord_x = 15;
defparam asyncreset_ctrl_X59_Y3_N0.coord_y = 12;
defparam asyncreset_ctrl_X59_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X59_Y3_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X59_Y4_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y4_SIG ));
defparam asyncreset_ctrl_X59_Y4_N0.coord_x = 17;
defparam asyncreset_ctrl_X59_Y4_N0.coord_y = 11;
defparam asyncreset_ctrl_X59_Y4_N0.coord_z = 0;
defparam asyncreset_ctrl_X59_Y4_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X59_Y5_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ));
defparam asyncreset_ctrl_X59_Y5_N0.coord_x = 14;
defparam asyncreset_ctrl_X59_Y5_N0.coord_y = 8;
defparam asyncreset_ctrl_X59_Y5_N0.coord_z = 0;
defparam asyncreset_ctrl_X59_Y5_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X59_Y6_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y6_SIG ));
defparam asyncreset_ctrl_X59_Y6_N0.coord_x = 18;
defparam asyncreset_ctrl_X59_Y6_N0.coord_y = 11;
defparam asyncreset_ctrl_X59_Y6_N0.coord_z = 0;
defparam asyncreset_ctrl_X59_Y6_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X59_Y7_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ));
defparam asyncreset_ctrl_X59_Y7_N0.coord_x = 18;
defparam asyncreset_ctrl_X59_Y7_N0.coord_y = 5;
defparam asyncreset_ctrl_X59_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X59_Y7_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X59_Y8_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ));
defparam asyncreset_ctrl_X59_Y8_N0.coord_x = 14;
defparam asyncreset_ctrl_X59_Y8_N0.coord_y = 6;
defparam asyncreset_ctrl_X59_Y8_N0.coord_z = 0;
defparam asyncreset_ctrl_X59_Y8_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X59_Y9_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ));
defparam asyncreset_ctrl_X59_Y9_N0.coord_x = 18;
defparam asyncreset_ctrl_X59_Y9_N0.coord_y = 10;
defparam asyncreset_ctrl_X59_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X59_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X60_Y10_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ));
defparam asyncreset_ctrl_X60_Y10_N0.coord_x = 20;
defparam asyncreset_ctrl_X60_Y10_N0.coord_y = 11;
defparam asyncreset_ctrl_X60_Y10_N0.coord_z = 0;
defparam asyncreset_ctrl_X60_Y10_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X60_Y11_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ));
defparam asyncreset_ctrl_X60_Y11_N0.coord_x = 19;
defparam asyncreset_ctrl_X60_Y11_N0.coord_y = 4;
defparam asyncreset_ctrl_X60_Y11_N0.coord_z = 0;
defparam asyncreset_ctrl_X60_Y11_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X60_Y12_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ));
defparam asyncreset_ctrl_X60_Y12_N0.coord_x = 20;
defparam asyncreset_ctrl_X60_Y12_N0.coord_y = 7;
defparam asyncreset_ctrl_X60_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X60_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X60_Y1_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ));
defparam asyncreset_ctrl_X60_Y1_N0.coord_x = 17;
defparam asyncreset_ctrl_X60_Y1_N0.coord_y = 1;
defparam asyncreset_ctrl_X60_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X60_Y1_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X60_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ));
defparam asyncreset_ctrl_X60_Y2_N0.coord_x = 11;
defparam asyncreset_ctrl_X60_Y2_N0.coord_y = 4;
defparam asyncreset_ctrl_X60_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X60_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X60_Y3_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y3_SIG ));
defparam asyncreset_ctrl_X60_Y3_N0.coord_x = 15;
defparam asyncreset_ctrl_X60_Y3_N0.coord_y = 7;
defparam asyncreset_ctrl_X60_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X60_Y3_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X60_Y4_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ));
defparam asyncreset_ctrl_X60_Y4_N0.coord_x = 15;
defparam asyncreset_ctrl_X60_Y4_N0.coord_y = 8;
defparam asyncreset_ctrl_X60_Y4_N0.coord_z = 0;
defparam asyncreset_ctrl_X60_Y4_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X60_Y5_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ));
defparam asyncreset_ctrl_X60_Y5_N0.coord_x = 15;
defparam asyncreset_ctrl_X60_Y5_N0.coord_y = 10;
defparam asyncreset_ctrl_X60_Y5_N0.coord_z = 0;
defparam asyncreset_ctrl_X60_Y5_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X60_Y6_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ));
defparam asyncreset_ctrl_X60_Y6_N0.coord_x = 18;
defparam asyncreset_ctrl_X60_Y6_N0.coord_y = 7;
defparam asyncreset_ctrl_X60_Y6_N0.coord_z = 0;
defparam asyncreset_ctrl_X60_Y6_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X60_Y7_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y7_SIG ));
defparam asyncreset_ctrl_X60_Y7_N0.coord_x = 18;
defparam asyncreset_ctrl_X60_Y7_N0.coord_y = 4;
defparam asyncreset_ctrl_X60_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X60_Y7_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X60_Y8_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ));
defparam asyncreset_ctrl_X60_Y8_N0.coord_x = 16;
defparam asyncreset_ctrl_X60_Y8_N0.coord_y = 7;
defparam asyncreset_ctrl_X60_Y8_N0.coord_z = 0;
defparam asyncreset_ctrl_X60_Y8_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X60_Y9_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ));
defparam asyncreset_ctrl_X60_Y9_N0.coord_x = 20;
defparam asyncreset_ctrl_X60_Y9_N0.coord_y = 4;
defparam asyncreset_ctrl_X60_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X60_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X61_Y10_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y10_SIG ));
defparam asyncreset_ctrl_X61_Y10_N0.coord_x = 19;
defparam asyncreset_ctrl_X61_Y10_N0.coord_y = 9;
defparam asyncreset_ctrl_X61_Y10_N0.coord_z = 0;
defparam asyncreset_ctrl_X61_Y10_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X61_Y11_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ));
defparam asyncreset_ctrl_X61_Y11_N0.coord_x = 19;
defparam asyncreset_ctrl_X61_Y11_N0.coord_y = 8;
defparam asyncreset_ctrl_X61_Y11_N0.coord_z = 0;
defparam asyncreset_ctrl_X61_Y11_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X61_Y12_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ));
defparam asyncreset_ctrl_X61_Y12_N0.coord_x = 19;
defparam asyncreset_ctrl_X61_Y12_N0.coord_y = 6;
defparam asyncreset_ctrl_X61_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X61_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X61_Y1_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ));
defparam asyncreset_ctrl_X61_Y1_N0.coord_x = 18;
defparam asyncreset_ctrl_X61_Y1_N0.coord_y = 1;
defparam asyncreset_ctrl_X61_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X61_Y1_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X61_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y2_SIG ));
defparam asyncreset_ctrl_X61_Y2_N0.coord_x = 15;
defparam asyncreset_ctrl_X61_Y2_N0.coord_y = 5;
defparam asyncreset_ctrl_X61_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X61_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X61_Y3_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ));
defparam asyncreset_ctrl_X61_Y3_N0.coord_x = 15;
defparam asyncreset_ctrl_X61_Y3_N0.coord_y = 1;
defparam asyncreset_ctrl_X61_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X61_Y3_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X61_Y4_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ));
defparam asyncreset_ctrl_X61_Y4_N0.coord_x = 17;
defparam asyncreset_ctrl_X61_Y4_N0.coord_y = 8;
defparam asyncreset_ctrl_X61_Y4_N0.coord_z = 0;
defparam asyncreset_ctrl_X61_Y4_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X61_Y5_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ));
defparam asyncreset_ctrl_X61_Y5_N0.coord_x = 14;
defparam asyncreset_ctrl_X61_Y5_N0.coord_y = 1;
defparam asyncreset_ctrl_X61_Y5_N0.coord_z = 0;
defparam asyncreset_ctrl_X61_Y5_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X61_Y6_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ));
defparam asyncreset_ctrl_X61_Y6_N0.coord_x = 15;
defparam asyncreset_ctrl_X61_Y6_N0.coord_y = 9;
defparam asyncreset_ctrl_X61_Y6_N0.coord_z = 0;
defparam asyncreset_ctrl_X61_Y6_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X61_Y7_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ));
defparam asyncreset_ctrl_X61_Y7_N0.coord_x = 17;
defparam asyncreset_ctrl_X61_Y7_N0.coord_y = 3;
defparam asyncreset_ctrl_X61_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X61_Y7_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X61_Y8_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ));
defparam asyncreset_ctrl_X61_Y8_N0.coord_x = 19;
defparam asyncreset_ctrl_X61_Y8_N0.coord_y = 2;
defparam asyncreset_ctrl_X61_Y8_N0.coord_z = 0;
defparam asyncreset_ctrl_X61_Y8_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X61_Y9_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ));
defparam asyncreset_ctrl_X61_Y9_N0.coord_x = 19;
defparam asyncreset_ctrl_X61_Y9_N0.coord_y = 7;
defparam asyncreset_ctrl_X61_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X61_Y9_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X62_Y10_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ));
defparam asyncreset_ctrl_X62_Y10_N0.coord_x = 20;
defparam asyncreset_ctrl_X62_Y10_N0.coord_y = 12;
defparam asyncreset_ctrl_X62_Y10_N0.coord_z = 0;
defparam asyncreset_ctrl_X62_Y10_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X62_Y11_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ));
defparam asyncreset_ctrl_X62_Y11_N0.coord_x = 20;
defparam asyncreset_ctrl_X62_Y11_N0.coord_y = 9;
defparam asyncreset_ctrl_X62_Y11_N0.coord_z = 0;
defparam asyncreset_ctrl_X62_Y11_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X62_Y12_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ));
defparam asyncreset_ctrl_X62_Y12_N0.coord_x = 20;
defparam asyncreset_ctrl_X62_Y12_N0.coord_y = 6;
defparam asyncreset_ctrl_X62_Y12_N0.coord_z = 0;
defparam asyncreset_ctrl_X62_Y12_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X62_Y1_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y1_SIG ));
defparam asyncreset_ctrl_X62_Y1_N0.coord_x = 12;
defparam asyncreset_ctrl_X62_Y1_N0.coord_y = 1;
defparam asyncreset_ctrl_X62_Y1_N0.coord_z = 0;
defparam asyncreset_ctrl_X62_Y1_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X62_Y2_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ));
defparam asyncreset_ctrl_X62_Y2_N0.coord_x = 17;
defparam asyncreset_ctrl_X62_Y2_N0.coord_y = 6;
defparam asyncreset_ctrl_X62_Y2_N0.coord_z = 0;
defparam asyncreset_ctrl_X62_Y2_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X62_Y3_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ));
defparam asyncreset_ctrl_X62_Y3_N0.coord_x = 16;
defparam asyncreset_ctrl_X62_Y3_N0.coord_y = 6;
defparam asyncreset_ctrl_X62_Y3_N0.coord_z = 0;
defparam asyncreset_ctrl_X62_Y3_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X62_Y4_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y4_SIG ));
defparam asyncreset_ctrl_X62_Y4_N0.coord_x = 14;
defparam asyncreset_ctrl_X62_Y4_N0.coord_y = 3;
defparam asyncreset_ctrl_X62_Y4_N0.coord_z = 0;
defparam asyncreset_ctrl_X62_Y4_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X62_Y5_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ));
defparam asyncreset_ctrl_X62_Y5_N0.coord_x = 17;
defparam asyncreset_ctrl_X62_Y5_N0.coord_y = 10;
defparam asyncreset_ctrl_X62_Y5_N0.coord_z = 0;
defparam asyncreset_ctrl_X62_Y5_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X62_Y6_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y6_SIG ));
defparam asyncreset_ctrl_X62_Y6_N0.coord_x = 17;
defparam asyncreset_ctrl_X62_Y6_N0.coord_y = 12;
defparam asyncreset_ctrl_X62_Y6_N0.coord_z = 0;
defparam asyncreset_ctrl_X62_Y6_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X62_Y7_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ));
defparam asyncreset_ctrl_X62_Y7_N0.coord_x = 15;
defparam asyncreset_ctrl_X62_Y7_N0.coord_y = 6;
defparam asyncreset_ctrl_X62_Y7_N0.coord_z = 0;
defparam asyncreset_ctrl_X62_Y7_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X62_Y8_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ));
defparam asyncreset_ctrl_X62_Y8_N0.coord_x = 18;
defparam asyncreset_ctrl_X62_Y8_N0.coord_y = 2;
defparam asyncreset_ctrl_X62_Y8_N0.coord_z = 0;
defparam asyncreset_ctrl_X62_Y8_N0.AsyncCtrlMux = 2'b10;

alta_asyncctrl asyncreset_ctrl_X62_Y9_N0(
	.Din(\sys_resetn~clkctrl_outclk ),
	.Dout(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ));
defparam asyncreset_ctrl_X62_Y9_N0.coord_x = 19;
defparam asyncreset_ctrl_X62_Y9_N0.coord_y = 11;
defparam asyncreset_ctrl_X62_Y9_N0.coord_z = 0;
defparam asyncreset_ctrl_X62_Y9_N0.AsyncCtrlMux = 2'b10;

alta_clkenctrl clken_ctrl_X43_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ));
defparam clken_ctrl_X43_Y2_N0.coord_x = 7;
defparam clken_ctrl_X43_Y2_N0.coord_y = 2;
defparam clken_ctrl_X43_Y2_N0.coord_z = 0;
defparam clken_ctrl_X43_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X43_Y2_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X46_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|load_counter[14]~19_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ));
defparam clken_ctrl_X46_Y2_N0.coord_x = 4;
defparam clken_ctrl_X46_Y2_N0.coord_y = 3;
defparam clken_ctrl_X46_Y2_N0.coord_z = 0;
defparam clken_ctrl_X46_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X46_Y2_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X46_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X46_Y3_SIG_VCC ));
defparam clken_ctrl_X46_Y3_N0.coord_x = 5;
defparam clken_ctrl_X46_Y3_N0.coord_y = 4;
defparam clken_ctrl_X46_Y3_N0.coord_z = 0;
defparam clken_ctrl_X46_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X46_Y3_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X47_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X47_Y2_SIG_VCC ));
defparam clken_ctrl_X47_Y2_N0.coord_x = 4;
defparam clken_ctrl_X47_Y2_N0.coord_y = 2;
defparam clken_ctrl_X47_Y2_N0.coord_z = 0;
defparam clken_ctrl_X47_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X47_Y2_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X47_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X47_Y3_SIG_VCC ));
defparam clken_ctrl_X47_Y3_N0.coord_x = 4;
defparam clken_ctrl_X47_Y3_N0.coord_y = 4;
defparam clken_ctrl_X47_Y3_N0.coord_z = 0;
defparam clken_ctrl_X47_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X47_Y3_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X48_Y1_N0(
	.ClkIn(\auto_generated_inst.hbo_13_1bc039b416d3bc4a_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_13_1bc039b416d3bc4a_bp_X48_Y1_SIG_VCC ));
defparam clken_ctrl_X48_Y1_N0.coord_x = 5;
defparam clken_ctrl_X48_Y1_N0.coord_y = 3;
defparam clken_ctrl_X48_Y1_N0.coord_z = 0;
defparam clken_ctrl_X48_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X48_Y1_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X48_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y2_SIG_VCC ));
defparam clken_ctrl_X48_Y2_N0.coord_x = 3;
defparam clken_ctrl_X48_Y2_N0.coord_y = 1;
defparam clken_ctrl_X48_Y2_N0.coord_z = 0;
defparam clken_ctrl_X48_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X48_Y2_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X48_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y3_SIG_VCC ));
defparam clken_ctrl_X48_Y3_N0.coord_x = 3;
defparam clken_ctrl_X48_Y3_N0.coord_y = 2;
defparam clken_ctrl_X48_Y3_N0.coord_z = 0;
defparam clken_ctrl_X48_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X48_Y3_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X49_Y1_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X49_Y1_SIG_VCC ));
defparam clken_ctrl_X49_Y1_N0.coord_x = 6;
defparam clken_ctrl_X49_Y1_N0.coord_y = 1;
defparam clken_ctrl_X49_Y1_N0.coord_z = 0;
defparam clken_ctrl_X49_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X49_Y1_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X49_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|capture_done~q ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X49_Y2_SIG_SIG ));
defparam clken_ctrl_X49_Y2_N0.coord_x = 9;
defparam clken_ctrl_X49_Y2_N0.coord_y = 3;
defparam clken_ctrl_X49_Y2_N0.coord_z = 0;
defparam clken_ctrl_X49_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X49_Y2_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X49_Y2_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|Decoder0~5_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~5_combout_X49_Y2_SIG_SIG ));
defparam clken_ctrl_X49_Y2_N1.coord_x = 9;
defparam clken_ctrl_X49_Y2_N1.coord_y = 3;
defparam clken_ctrl_X49_Y2_N1.coord_z = 1;
defparam clken_ctrl_X49_Y2_N1.ClkMux = 2'b10;
defparam clken_ctrl_X49_Y2_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X49_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|Decoder0~4_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~4_combout_X49_Y3_SIG_SIG ));
defparam clken_ctrl_X49_Y3_N0.coord_x = 6;
defparam clken_ctrl_X49_Y3_N0.coord_y = 4;
defparam clken_ctrl_X49_Y3_N0.coord_z = 0;
defparam clken_ctrl_X49_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X49_Y3_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X49_Y3_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|Decoder0~7_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~7_combout_X49_Y3_SIG_SIG ));
defparam clken_ctrl_X49_Y3_N1.coord_x = 6;
defparam clken_ctrl_X49_Y3_N1.coord_y = 4;
defparam clken_ctrl_X49_Y3_N1.coord_z = 1;
defparam clken_ctrl_X49_Y3_N1.ClkMux = 2'b10;
defparam clken_ctrl_X49_Y3_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X49_Y4_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|capture_done~q ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X49_Y4_SIG_SIG ));
defparam clken_ctrl_X49_Y4_N0.coord_x = 3;
defparam clken_ctrl_X49_Y4_N0.coord_y = 4;
defparam clken_ctrl_X49_Y4_N0.coord_z = 0;
defparam clken_ctrl_X49_Y4_N0.ClkMux = 2'b10;
defparam clken_ctrl_X49_Y4_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X49_Y4_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X49_Y4_SIG_VCC ));
defparam clken_ctrl_X49_Y4_N1.coord_x = 3;
defparam clken_ctrl_X49_Y4_N1.coord_y = 4;
defparam clken_ctrl_X49_Y4_N1.coord_z = 1;
defparam clken_ctrl_X49_Y4_N1.ClkMux = 2'b10;
defparam clken_ctrl_X49_Y4_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X50_Y1_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|Equal0~0_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|Equal0~0_combout_X50_Y1_SIG_INV ));
defparam clken_ctrl_X50_Y1_N0.coord_x = 7;
defparam clken_ctrl_X50_Y1_N0.coord_y = 1;
defparam clken_ctrl_X50_Y1_N0.coord_z = 0;
defparam clken_ctrl_X50_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X50_Y1_N0.ClkEnMux = 2'b11;

alta_clkenctrl clken_ctrl_X50_Y1_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X50_Y1_SIG_VCC ));
defparam clken_ctrl_X50_Y1_N1.coord_x = 7;
defparam clken_ctrl_X50_Y1_N1.coord_y = 1;
defparam clken_ctrl_X50_Y1_N1.coord_z = 1;
defparam clken_ctrl_X50_Y1_N1.ClkMux = 2'b10;
defparam clken_ctrl_X50_Y1_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X50_Y2_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|bit_counter[7]~8_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|bit_counter[7]~8_combout_X50_Y2_SIG_SIG ));
defparam clken_ctrl_X50_Y2_N1.coord_x = 9;
defparam clken_ctrl_X50_Y2_N1.coord_y = 2;
defparam clken_ctrl_X50_Y2_N1.coord_z = 1;
defparam clken_ctrl_X50_Y2_N1.ClkMux = 2'b10;
defparam clken_ctrl_X50_Y2_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X50_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|Decoder0~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~1_combout_X50_Y3_SIG_SIG ));
defparam clken_ctrl_X50_Y3_N0.coord_x = 8;
defparam clken_ctrl_X50_Y3_N0.coord_y = 4;
defparam clken_ctrl_X50_Y3_N0.coord_z = 0;
defparam clken_ctrl_X50_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X50_Y3_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X50_Y3_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|Decoder0~8_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~8_combout_X50_Y3_SIG_SIG ));
defparam clken_ctrl_X50_Y3_N1.coord_x = 8;
defparam clken_ctrl_X50_Y3_N1.coord_y = 4;
defparam clken_ctrl_X50_Y3_N1.coord_z = 1;
defparam clken_ctrl_X50_Y3_N1.ClkMux = 2'b10;
defparam clken_ctrl_X50_Y3_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X50_Y4_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X50_Y4_SIG_SIG ));
defparam clken_ctrl_X50_Y4_N0.coord_x = 9;
defparam clken_ctrl_X50_Y4_N0.coord_y = 1;
defparam clken_ctrl_X50_Y4_N0.coord_z = 0;
defparam clken_ctrl_X50_Y4_N0.ClkMux = 2'b10;
defparam clken_ctrl_X50_Y4_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X51_Y1_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|scaler_counter[0]~0_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|scaler_counter[0]~0_combout_X51_Y1_SIG_SIG ));
defparam clken_ctrl_X51_Y1_N0.coord_x = 8;
defparam clken_ctrl_X51_Y1_N0.coord_y = 1;
defparam clken_ctrl_X51_Y1_N0.coord_z = 0;
defparam clken_ctrl_X51_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X51_Y1_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X51_Y1_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X51_Y1_SIG_VCC ));
defparam clken_ctrl_X51_Y1_N1.coord_x = 8;
defparam clken_ctrl_X51_Y1_N1.coord_y = 1;
defparam clken_ctrl_X51_Y1_N1.coord_z = 1;
defparam clken_ctrl_X51_Y1_N1.ClkMux = 2'b10;
defparam clken_ctrl_X51_Y1_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X51_Y2_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|byte_counter[4]~10_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|byte_counter[4]~10_combout_X51_Y2_SIG_SIG ));
defparam clken_ctrl_X51_Y2_N1.coord_x = 8;
defparam clken_ctrl_X51_Y2_N1.coord_y = 2;
defparam clken_ctrl_X51_Y2_N1.coord_z = 1;
defparam clken_ctrl_X51_Y2_N1.ClkMux = 2'b10;
defparam clken_ctrl_X51_Y2_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X51_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|Decoder0~2_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~2_combout_X51_Y3_SIG_SIG ));
defparam clken_ctrl_X51_Y3_N0.coord_x = 9;
defparam clken_ctrl_X51_Y3_N0.coord_y = 4;
defparam clken_ctrl_X51_Y3_N0.coord_z = 0;
defparam clken_ctrl_X51_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X51_Y3_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X51_Y3_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|capture_done~q ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X51_Y3_SIG_SIG ));
defparam clken_ctrl_X51_Y3_N1.coord_x = 9;
defparam clken_ctrl_X51_Y3_N1.coord_y = 4;
defparam clken_ctrl_X51_Y3_N1.coord_z = 1;
defparam clken_ctrl_X51_Y3_N1.ClkMux = 2'b10;
defparam clken_ctrl_X51_Y3_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X51_Y4_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ));
defparam clken_ctrl_X51_Y4_N0.coord_x = 15;
defparam clken_ctrl_X51_Y4_N0.coord_y = 2;
defparam clken_ctrl_X51_Y4_N0.coord_z = 0;
defparam clken_ctrl_X51_Y4_N0.ClkMux = 2'b10;
defparam clken_ctrl_X51_Y4_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X51_Y4_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|sdata_reg[0]~0_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X51_Y4_SIG_SIG ));
defparam clken_ctrl_X51_Y4_N1.coord_x = 15;
defparam clken_ctrl_X51_Y4_N1.coord_y = 2;
defparam clken_ctrl_X51_Y4_N1.coord_z = 1;
defparam clken_ctrl_X51_Y4_N1.ClkMux = 2'b10;
defparam clken_ctrl_X51_Y4_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X52_Y1_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ));
defparam clken_ctrl_X52_Y1_N0.coord_x = 11;
defparam clken_ctrl_X52_Y1_N0.coord_y = 1;
defparam clken_ctrl_X52_Y1_N0.coord_z = 0;
defparam clken_ctrl_X52_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X52_Y1_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X52_Y1_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|sdata_reg[0]~0_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X52_Y1_SIG_SIG ));
defparam clken_ctrl_X52_Y1_N1.coord_x = 11;
defparam clken_ctrl_X52_Y1_N1.coord_y = 1;
defparam clken_ctrl_X52_Y1_N1.coord_z = 1;
defparam clken_ctrl_X52_Y1_N1.ClkMux = 2'b10;
defparam clken_ctrl_X52_Y1_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X52_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|sdata_reg[0]~0_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X52_Y2_SIG_SIG ));
defparam clken_ctrl_X52_Y2_N0.coord_x = 16;
defparam clken_ctrl_X52_Y2_N0.coord_y = 5;
defparam clken_ctrl_X52_Y2_N0.coord_z = 0;
defparam clken_ctrl_X52_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X52_Y2_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X52_Y2_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ));
defparam clken_ctrl_X52_Y2_N1.coord_x = 16;
defparam clken_ctrl_X52_Y2_N1.coord_y = 5;
defparam clken_ctrl_X52_Y2_N1.coord_z = 1;
defparam clken_ctrl_X52_Y2_N1.ClkMux = 2'b10;
defparam clken_ctrl_X52_Y2_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X52_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|Decoder0~3_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~3_combout_X52_Y3_SIG_SIG ));
defparam clken_ctrl_X52_Y3_N0.coord_x = 8;
defparam clken_ctrl_X52_Y3_N0.coord_y = 3;
defparam clken_ctrl_X52_Y3_N0.coord_z = 0;
defparam clken_ctrl_X52_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X52_Y3_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X52_Y3_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|Decoder0~6_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~6_combout_X52_Y3_SIG_SIG ));
defparam clken_ctrl_X52_Y3_N1.coord_x = 8;
defparam clken_ctrl_X52_Y3_N1.coord_y = 3;
defparam clken_ctrl_X52_Y3_N1.coord_z = 1;
defparam clken_ctrl_X52_Y3_N1.ClkMux = 2'b10;
defparam clken_ctrl_X52_Y3_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X52_Y4_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ));
defparam clken_ctrl_X52_Y4_N0.coord_x = 16;
defparam clken_ctrl_X52_Y4_N0.coord_y = 2;
defparam clken_ctrl_X52_Y4_N0.coord_z = 0;
defparam clken_ctrl_X52_Y4_N0.ClkMux = 2'b10;
defparam clken_ctrl_X52_Y4_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X53_Y1_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ));
defparam clken_ctrl_X53_Y1_N0.coord_x = 16;
defparam clken_ctrl_X53_Y1_N0.coord_y = 1;
defparam clken_ctrl_X53_Y1_N0.coord_z = 0;
defparam clken_ctrl_X53_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X53_Y1_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X53_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ));
defparam clken_ctrl_X53_Y2_N0.coord_x = 19;
defparam clken_ctrl_X53_Y2_N0.coord_y = 5;
defparam clken_ctrl_X53_Y2_N0.coord_z = 0;
defparam clken_ctrl_X53_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X53_Y2_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X53_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|capture_done~q ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ));
defparam clken_ctrl_X53_Y3_N0.coord_x = 7;
defparam clken_ctrl_X53_Y3_N0.coord_y = 4;
defparam clken_ctrl_X53_Y3_N0.coord_z = 0;
defparam clken_ctrl_X53_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X53_Y3_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X53_Y4_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ));
defparam clken_ctrl_X53_Y4_N0.coord_x = 15;
defparam clken_ctrl_X53_Y4_N0.coord_y = 4;
defparam clken_ctrl_X53_Y4_N0.coord_z = 0;
defparam clken_ctrl_X53_Y4_N0.ClkMux = 2'b10;
defparam clken_ctrl_X53_Y4_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X53_Y4_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|sdata_reg[0]~0_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X53_Y4_SIG_SIG ));
defparam clken_ctrl_X53_Y4_N1.coord_x = 15;
defparam clken_ctrl_X53_Y4_N1.coord_y = 4;
defparam clken_ctrl_X53_Y4_N1.coord_z = 1;
defparam clken_ctrl_X53_Y4_N1.ClkMux = 2'b10;
defparam clken_ctrl_X53_Y4_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X54_Y1_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|sdata_reg[0]~0_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ));
defparam clken_ctrl_X54_Y1_N0.coord_x = 20;
defparam clken_ctrl_X54_Y1_N0.coord_y = 2;
defparam clken_ctrl_X54_Y1_N0.coord_z = 0;
defparam clken_ctrl_X54_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X54_Y1_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X54_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X54_Y2_SIG_VCC ));
defparam clken_ctrl_X54_Y2_N0.coord_x = 14;
defparam clken_ctrl_X54_Y2_N0.coord_y = 5;
defparam clken_ctrl_X54_Y2_N0.coord_z = 0;
defparam clken_ctrl_X54_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X54_Y2_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X54_Y2_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~52_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X54_Y2_SIG_SIG ));
defparam clken_ctrl_X54_Y2_N1.coord_x = 14;
defparam clken_ctrl_X54_Y2_N1.coord_y = 5;
defparam clken_ctrl_X54_Y2_N1.coord_z = 1;
defparam clken_ctrl_X54_Y2_N1.ClkMux = 2'b10;
defparam clken_ctrl_X54_Y2_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X54_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|ahb_read_transfer~combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X54_Y3_SIG_SIG ));
defparam clken_ctrl_X54_Y3_N0.coord_x = 14;
defparam clken_ctrl_X54_Y3_N0.coord_y = 12;
defparam clken_ctrl_X54_Y3_N0.coord_z = 0;
defparam clken_ctrl_X54_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X54_Y3_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X54_Y3_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|Equal2~0_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X54_Y3_SIG_SIG ));
defparam clken_ctrl_X54_Y3_N1.coord_x = 14;
defparam clken_ctrl_X54_Y3_N1.coord_y = 12;
defparam clken_ctrl_X54_Y3_N1.coord_z = 1;
defparam clken_ctrl_X54_Y3_N1.ClkMux = 2'b10;
defparam clken_ctrl_X54_Y3_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X54_Y4_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~79_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X54_Y4_SIG_SIG ));
defparam clken_ctrl_X54_Y4_N0.coord_x = 11;
defparam clken_ctrl_X54_Y4_N0.coord_y = 2;
defparam clken_ctrl_X54_Y4_N0.coord_z = 0;
defparam clken_ctrl_X54_Y4_N0.ClkMux = 2'b10;
defparam clken_ctrl_X54_Y4_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X54_Y4_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X54_Y4_SIG_VCC ));
defparam clken_ctrl_X54_Y4_N1.coord_x = 11;
defparam clken_ctrl_X54_Y4_N1.coord_y = 2;
defparam clken_ctrl_X54_Y4_N1.coord_z = 1;
defparam clken_ctrl_X54_Y4_N1.ClkMux = 2'b10;
defparam clken_ctrl_X54_Y4_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X56_Y10_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y10_SIG_VCC ));
defparam clken_ctrl_X56_Y10_N0.coord_x = 11;
defparam clken_ctrl_X56_Y10_N0.coord_y = 3;
defparam clken_ctrl_X56_Y10_N0.coord_z = 0;
defparam clken_ctrl_X56_Y10_N0.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y10_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X56_Y10_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~50_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X56_Y10_SIG_SIG ));
defparam clken_ctrl_X56_Y10_N1.coord_x = 11;
defparam clken_ctrl_X56_Y10_N1.coord_y = 3;
defparam clken_ctrl_X56_Y10_N1.coord_z = 1;
defparam clken_ctrl_X56_Y10_N1.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y10_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y11_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y11_SIG_SIG ));
defparam clken_ctrl_X56_Y11_N0.coord_x = 19;
defparam clken_ctrl_X56_Y11_N0.coord_y = 10;
defparam clken_ctrl_X56_Y11_N0.coord_z = 0;
defparam clken_ctrl_X56_Y11_N0.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y11_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y11_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y11_SIG_VCC ));
defparam clken_ctrl_X56_Y11_N1.coord_x = 19;
defparam clken_ctrl_X56_Y11_N1.coord_y = 10;
defparam clken_ctrl_X56_Y11_N1.coord_z = 1;
defparam clken_ctrl_X56_Y11_N1.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y11_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X56_Y12_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ));
defparam clken_ctrl_X56_Y12_N0.coord_x = 20;
defparam clken_ctrl_X56_Y12_N0.coord_y = 8;
defparam clken_ctrl_X56_Y12_N0.coord_z = 0;
defparam clken_ctrl_X56_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y12_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y1_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~54_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X56_Y1_SIG_SIG ));
defparam clken_ctrl_X56_Y1_N0.coord_x = 10;
defparam clken_ctrl_X56_Y1_N0.coord_y = 2;
defparam clken_ctrl_X56_Y1_N0.coord_z = 0;
defparam clken_ctrl_X56_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y1_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y1_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y1_SIG_VCC ));
defparam clken_ctrl_X56_Y1_N1.coord_x = 10;
defparam clken_ctrl_X56_Y1_N1.coord_y = 2;
defparam clken_ctrl_X56_Y1_N1.coord_z = 1;
defparam clken_ctrl_X56_Y1_N1.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y1_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X56_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~78_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X56_Y2_SIG_SIG ));
defparam clken_ctrl_X56_Y2_N0.coord_x = 16;
defparam clken_ctrl_X56_Y2_N0.coord_y = 11;
defparam clken_ctrl_X56_Y2_N0.coord_z = 0;
defparam clken_ctrl_X56_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y2_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y2_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~17_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X56_Y2_SIG_SIG ));
defparam clken_ctrl_X56_Y2_N1.coord_x = 16;
defparam clken_ctrl_X56_Y2_N1.coord_y = 11;
defparam clken_ctrl_X56_Y2_N1.coord_z = 1;
defparam clken_ctrl_X56_Y2_N1.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y2_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|ahb_read_transfer~combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y3_SIG_SIG ));
defparam clken_ctrl_X56_Y3_N0.coord_x = 12;
defparam clken_ctrl_X56_Y3_N0.coord_y = 4;
defparam clken_ctrl_X56_Y3_N0.coord_z = 0;
defparam clken_ctrl_X56_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y3_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y3_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|capture_done~q ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y3_SIG_SIG ));
defparam clken_ctrl_X56_Y3_N1.coord_x = 12;
defparam clken_ctrl_X56_Y3_N1.coord_y = 4;
defparam clken_ctrl_X56_Y3_N1.coord_z = 1;
defparam clken_ctrl_X56_Y3_N1.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y3_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y4_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y4_SIG_VCC ));
defparam clken_ctrl_X56_Y4_N0.coord_x = 17;
defparam clken_ctrl_X56_Y4_N0.coord_y = 4;
defparam clken_ctrl_X56_Y4_N0.coord_z = 0;
defparam clken_ctrl_X56_Y4_N0.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y4_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X56_Y4_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~61_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X56_Y4_SIG_SIG ));
defparam clken_ctrl_X56_Y4_N1.coord_x = 17;
defparam clken_ctrl_X56_Y4_N1.coord_y = 4;
defparam clken_ctrl_X56_Y4_N1.coord_z = 1;
defparam clken_ctrl_X56_Y4_N1.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y4_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y5_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|capture_done~q ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y5_SIG_SIG ));
defparam clken_ctrl_X56_Y5_N0.coord_x = 10;
defparam clken_ctrl_X56_Y5_N0.coord_y = 4;
defparam clken_ctrl_X56_Y5_N0.coord_z = 0;
defparam clken_ctrl_X56_Y5_N0.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y5_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y5_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|ahb_read_transfer~combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y5_SIG_SIG ));
defparam clken_ctrl_X56_Y5_N1.coord_x = 10;
defparam clken_ctrl_X56_Y5_N1.coord_y = 4;
defparam clken_ctrl_X56_Y5_N1.coord_z = 1;
defparam clken_ctrl_X56_Y5_N1.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y5_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y6_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y6_SIG_VCC ));
defparam clken_ctrl_X56_Y6_N0.coord_x = 17;
defparam clken_ctrl_X56_Y6_N0.coord_y = 2;
defparam clken_ctrl_X56_Y6_N0.coord_z = 0;
defparam clken_ctrl_X56_Y6_N0.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y6_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X56_Y6_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~57_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X56_Y6_SIG_SIG ));
defparam clken_ctrl_X56_Y6_N1.coord_x = 17;
defparam clken_ctrl_X56_Y6_N1.coord_y = 2;
defparam clken_ctrl_X56_Y6_N1.coord_z = 1;
defparam clken_ctrl_X56_Y6_N1.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y6_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y7_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~58_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y7_SIG_SIG ));
defparam clken_ctrl_X56_Y7_N0.coord_x = 14;
defparam clken_ctrl_X56_Y7_N0.coord_y = 2;
defparam clken_ctrl_X56_Y7_N0.coord_z = 0;
defparam clken_ctrl_X56_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y7_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y7_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y7_SIG_VCC ));
defparam clken_ctrl_X56_Y7_N1.coord_x = 14;
defparam clken_ctrl_X56_Y7_N1.coord_y = 2;
defparam clken_ctrl_X56_Y7_N1.coord_z = 1;
defparam clken_ctrl_X56_Y7_N1.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y7_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X56_Y8_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~33_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X56_Y8_SIG_SIG ));
defparam clken_ctrl_X56_Y8_N0.coord_x = 19;
defparam clken_ctrl_X56_Y8_N0.coord_y = 1;
defparam clken_ctrl_X56_Y8_N0.coord_z = 0;
defparam clken_ctrl_X56_Y8_N0.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y8_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y8_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~58_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y8_SIG_SIG ));
defparam clken_ctrl_X56_Y8_N1.coord_x = 19;
defparam clken_ctrl_X56_Y8_N1.coord_y = 1;
defparam clken_ctrl_X56_Y8_N1.coord_z = 1;
defparam clken_ctrl_X56_Y8_N1.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y8_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X56_Y9_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y9_SIG_VCC ));
defparam clken_ctrl_X56_Y9_N0.coord_x = 17;
defparam clken_ctrl_X56_Y9_N0.coord_y = 9;
defparam clken_ctrl_X56_Y9_N0.coord_z = 0;
defparam clken_ctrl_X56_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y9_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X56_Y9_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~56_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X56_Y9_SIG_SIG ));
defparam clken_ctrl_X56_Y9_N1.coord_x = 17;
defparam clken_ctrl_X56_Y9_N1.coord_y = 9;
defparam clken_ctrl_X56_Y9_N1.coord_z = 1;
defparam clken_ctrl_X56_Y9_N1.ClkMux = 2'b10;
defparam clken_ctrl_X56_Y9_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y10_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~65_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y10_SIG_SIG ));
defparam clken_ctrl_X57_Y10_N0.coord_x = 12;
defparam clken_ctrl_X57_Y10_N0.coord_y = 3;
defparam clken_ctrl_X57_Y10_N0.coord_z = 0;
defparam clken_ctrl_X57_Y10_N0.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y10_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y10_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~50_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X57_Y10_SIG_SIG ));
defparam clken_ctrl_X57_Y10_N1.coord_x = 12;
defparam clken_ctrl_X57_Y10_N1.coord_y = 3;
defparam clken_ctrl_X57_Y10_N1.coord_z = 1;
defparam clken_ctrl_X57_Y10_N1.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y10_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y11_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~25_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X57_Y11_SIG_SIG ));
defparam clken_ctrl_X57_Y11_N0.coord_x = 20;
defparam clken_ctrl_X57_Y11_N0.coord_y = 10;
defparam clken_ctrl_X57_Y11_N0.coord_z = 0;
defparam clken_ctrl_X57_Y11_N0.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y11_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y11_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~76_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X57_Y11_SIG_SIG ));
defparam clken_ctrl_X57_Y11_N1.coord_x = 20;
defparam clken_ctrl_X57_Y11_N1.coord_y = 10;
defparam clken_ctrl_X57_Y11_N1.coord_z = 1;
defparam clken_ctrl_X57_Y11_N1.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y11_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y12_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y12_SIG_VCC ));
defparam clken_ctrl_X57_Y12_N0.coord_x = 18;
defparam clken_ctrl_X57_Y12_N0.coord_y = 8;
defparam clken_ctrl_X57_Y12_N0.coord_z = 0;
defparam clken_ctrl_X57_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y12_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X57_Y12_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~65_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y12_SIG_SIG ));
defparam clken_ctrl_X57_Y12_N1.coord_x = 18;
defparam clken_ctrl_X57_Y12_N1.coord_y = 8;
defparam clken_ctrl_X57_Y12_N1.coord_z = 1;
defparam clken_ctrl_X57_Y12_N1.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y12_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y1_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y1_SIG_VCC ));
defparam clken_ctrl_X57_Y1_N0.coord_x = 12;
defparam clken_ctrl_X57_Y1_N0.coord_y = 2;
defparam clken_ctrl_X57_Y1_N0.coord_z = 0;
defparam clken_ctrl_X57_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y1_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X57_Y1_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~70_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X57_Y1_SIG_SIG ));
defparam clken_ctrl_X57_Y1_N1.coord_x = 12;
defparam clken_ctrl_X57_Y1_N1.coord_y = 2;
defparam clken_ctrl_X57_Y1_N1.coord_z = 1;
defparam clken_ctrl_X57_Y1_N1.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y1_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~17_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X57_Y2_SIG_SIG ));
defparam clken_ctrl_X57_Y2_N0.coord_x = 18;
defparam clken_ctrl_X57_Y2_N0.coord_y = 12;
defparam clken_ctrl_X57_Y2_N0.coord_z = 0;
defparam clken_ctrl_X57_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y2_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y2_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y2_SIG_VCC ));
defparam clken_ctrl_X57_Y2_N1.coord_x = 18;
defparam clken_ctrl_X57_Y2_N1.coord_y = 12;
defparam clken_ctrl_X57_Y2_N1.coord_z = 1;
defparam clken_ctrl_X57_Y2_N1.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y2_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X57_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|Equal2~0_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X57_Y3_SIG_SIG ));
defparam clken_ctrl_X57_Y3_N0.coord_x = 14;
defparam clken_ctrl_X57_Y3_N0.coord_y = 11;
defparam clken_ctrl_X57_Y3_N0.coord_z = 0;
defparam clken_ctrl_X57_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y3_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y3_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y3_SIG_VCC ));
defparam clken_ctrl_X57_Y3_N1.coord_x = 14;
defparam clken_ctrl_X57_Y3_N1.coord_y = 11;
defparam clken_ctrl_X57_Y3_N1.coord_z = 1;
defparam clken_ctrl_X57_Y3_N1.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y3_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X57_Y4_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y4_SIG_VCC ));
defparam clken_ctrl_X57_Y4_N0.coord_x = 16;
defparam clken_ctrl_X57_Y4_N0.coord_y = 4;
defparam clken_ctrl_X57_Y4_N0.coord_z = 0;
defparam clken_ctrl_X57_Y4_N0.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y4_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X57_Y4_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~30_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X57_Y4_SIG_SIG ));
defparam clken_ctrl_X57_Y4_N1.coord_x = 16;
defparam clken_ctrl_X57_Y4_N1.coord_y = 4;
defparam clken_ctrl_X57_Y4_N1.coord_z = 1;
defparam clken_ctrl_X57_Y4_N1.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y4_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y5_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|serial_lim_input_inst|ahb_read_transfer~combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X57_Y5_SIG_SIG ));
defparam clken_ctrl_X57_Y5_N1.coord_x = 14;
defparam clken_ctrl_X57_Y5_N1.coord_y = 7;
defparam clken_ctrl_X57_Y5_N1.coord_z = 1;
defparam clken_ctrl_X57_Y5_N1.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y5_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y6_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~14_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X57_Y6_SIG_SIG ));
defparam clken_ctrl_X57_Y6_N0.coord_x = 14;
defparam clken_ctrl_X57_Y6_N0.coord_y = 10;
defparam clken_ctrl_X57_Y6_N0.coord_z = 0;
defparam clken_ctrl_X57_Y6_N0.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y6_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y6_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~39_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X57_Y6_SIG_SIG ));
defparam clken_ctrl_X57_Y6_N1.coord_x = 14;
defparam clken_ctrl_X57_Y6_N1.coord_y = 10;
defparam clken_ctrl_X57_Y6_N1.coord_z = 1;
defparam clken_ctrl_X57_Y6_N1.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y6_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y7_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y7_SIG_VCC ));
defparam clken_ctrl_X57_Y7_N0.coord_x = 15;
defparam clken_ctrl_X57_Y7_N0.coord_y = 3;
defparam clken_ctrl_X57_Y7_N0.coord_z = 0;
defparam clken_ctrl_X57_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y7_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X57_Y7_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~39_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X57_Y7_SIG_SIG ));
defparam clken_ctrl_X57_Y7_N1.coord_x = 15;
defparam clken_ctrl_X57_Y7_N1.coord_y = 3;
defparam clken_ctrl_X57_Y7_N1.coord_z = 1;
defparam clken_ctrl_X57_Y7_N1.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y7_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y8_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~23_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X57_Y8_SIG_SIG ));
defparam clken_ctrl_X57_Y8_N0.coord_x = 18;
defparam clken_ctrl_X57_Y8_N0.coord_y = 3;
defparam clken_ctrl_X57_Y8_N0.coord_z = 0;
defparam clken_ctrl_X57_Y8_N0.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y8_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y8_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~62_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X57_Y8_SIG_SIG ));
defparam clken_ctrl_X57_Y8_N1.coord_x = 18;
defparam clken_ctrl_X57_Y8_N1.coord_y = 3;
defparam clken_ctrl_X57_Y8_N1.coord_z = 1;
defparam clken_ctrl_X57_Y8_N1.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y8_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y9_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~59_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X57_Y9_SIG_SIG ));
defparam clken_ctrl_X57_Y9_N0.coord_x = 16;
defparam clken_ctrl_X57_Y9_N0.coord_y = 9;
defparam clken_ctrl_X57_Y9_N0.coord_z = 0;
defparam clken_ctrl_X57_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y9_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X57_Y9_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y9_SIG_VCC ));
defparam clken_ctrl_X57_Y9_N1.coord_x = 16;
defparam clken_ctrl_X57_Y9_N1.coord_y = 9;
defparam clken_ctrl_X57_Y9_N1.coord_z = 1;
defparam clken_ctrl_X57_Y9_N1.ClkMux = 2'b10;
defparam clken_ctrl_X57_Y9_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X58_Y10_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~39_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X58_Y10_SIG_SIG ));
defparam clken_ctrl_X58_Y10_N0.coord_x = 17;
defparam clken_ctrl_X58_Y10_N0.coord_y = 7;
defparam clken_ctrl_X58_Y10_N0.coord_z = 0;
defparam clken_ctrl_X58_Y10_N0.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y10_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y10_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~42_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X58_Y10_SIG_SIG ));
defparam clken_ctrl_X58_Y10_N1.coord_x = 17;
defparam clken_ctrl_X58_Y10_N1.coord_y = 7;
defparam clken_ctrl_X58_Y10_N1.coord_z = 1;
defparam clken_ctrl_X58_Y10_N1.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y10_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y11_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~76_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X58_Y11_SIG_SIG ));
defparam clken_ctrl_X58_Y11_N0.coord_x = 19;
defparam clken_ctrl_X58_Y11_N0.coord_y = 12;
defparam clken_ctrl_X58_Y11_N0.coord_z = 0;
defparam clken_ctrl_X58_Y11_N0.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y11_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y11_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y11_SIG_VCC ));
defparam clken_ctrl_X58_Y11_N1.coord_x = 19;
defparam clken_ctrl_X58_Y11_N1.coord_y = 12;
defparam clken_ctrl_X58_Y11_N1.coord_z = 1;
defparam clken_ctrl_X58_Y11_N1.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y11_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X58_Y12_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y12_SIG_VCC ));
defparam clken_ctrl_X58_Y12_N0.coord_x = 20;
defparam clken_ctrl_X58_Y12_N0.coord_y = 3;
defparam clken_ctrl_X58_Y12_N0.coord_z = 0;
defparam clken_ctrl_X58_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y12_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X58_Y12_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~43_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X58_Y12_SIG_SIG ));
defparam clken_ctrl_X58_Y12_N1.coord_x = 20;
defparam clken_ctrl_X58_Y12_N1.coord_y = 3;
defparam clken_ctrl_X58_Y12_N1.coord_z = 1;
defparam clken_ctrl_X58_Y12_N1.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y12_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y1_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~70_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X58_Y1_SIG_SIG ));
defparam clken_ctrl_X58_Y1_N0.coord_x = 10;
defparam clken_ctrl_X58_Y1_N0.coord_y = 1;
defparam clken_ctrl_X58_Y1_N0.coord_z = 0;
defparam clken_ctrl_X58_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y1_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y1_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~54_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X58_Y1_SIG_SIG ));
defparam clken_ctrl_X58_Y1_N1.coord_x = 10;
defparam clken_ctrl_X58_Y1_N1.coord_y = 1;
defparam clken_ctrl_X58_Y1_N1.coord_z = 1;
defparam clken_ctrl_X58_Y1_N1.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y1_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~72_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X58_Y2_SIG_SIG ));
defparam clken_ctrl_X58_Y2_N0.coord_x = 16;
defparam clken_ctrl_X58_Y2_N0.coord_y = 10;
defparam clken_ctrl_X58_Y2_N0.coord_z = 0;
defparam clken_ctrl_X58_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y2_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y2_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~30_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X58_Y2_SIG_SIG ));
defparam clken_ctrl_X58_Y2_N1.coord_x = 16;
defparam clken_ctrl_X58_Y2_N1.coord_y = 10;
defparam clken_ctrl_X58_Y2_N1.coord_z = 1;
defparam clken_ctrl_X58_Y2_N1.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y2_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|Equal2~0_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X58_Y3_SIG_SIG ));
defparam clken_ctrl_X58_Y3_N0.coord_x = 15;
defparam clken_ctrl_X58_Y3_N0.coord_y = 11;
defparam clken_ctrl_X58_Y3_N0.coord_z = 0;
defparam clken_ctrl_X58_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y3_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y3_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~14_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X58_Y3_SIG_SIG ));
defparam clken_ctrl_X58_Y3_N1.coord_x = 15;
defparam clken_ctrl_X58_Y3_N1.coord_y = 11;
defparam clken_ctrl_X58_Y3_N1.coord_z = 1;
defparam clken_ctrl_X58_Y3_N1.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y3_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y4_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~45_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X58_Y4_SIG_SIG ));
defparam clken_ctrl_X58_Y4_N0.coord_x = 16;
defparam clken_ctrl_X58_Y4_N0.coord_y = 8;
defparam clken_ctrl_X58_Y4_N0.coord_z = 0;
defparam clken_ctrl_X58_Y4_N0.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y4_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y4_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y4_SIG_VCC ));
defparam clken_ctrl_X58_Y4_N1.coord_x = 16;
defparam clken_ctrl_X58_Y4_N1.coord_y = 8;
defparam clken_ctrl_X58_Y4_N1.coord_z = 1;
defparam clken_ctrl_X58_Y4_N1.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y4_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X58_Y5_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~24_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X58_Y5_SIG_SIG ));
defparam clken_ctrl_X58_Y5_N0.coord_x = 16;
defparam clken_ctrl_X58_Y5_N0.coord_y = 12;
defparam clken_ctrl_X58_Y5_N0.coord_z = 0;
defparam clken_ctrl_X58_Y5_N0.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y5_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y5_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~14_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X58_Y5_SIG_SIG ));
defparam clken_ctrl_X58_Y5_N1.coord_x = 16;
defparam clken_ctrl_X58_Y5_N1.coord_y = 12;
defparam clken_ctrl_X58_Y5_N1.coord_z = 1;
defparam clken_ctrl_X58_Y5_N1.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y5_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y6_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~44_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X58_Y6_SIG_SIG ));
defparam clken_ctrl_X58_Y6_N0.coord_x = 14;
defparam clken_ctrl_X58_Y6_N0.coord_y = 9;
defparam clken_ctrl_X58_Y6_N0.coord_z = 0;
defparam clken_ctrl_X58_Y6_N0.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y6_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y6_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~79_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X58_Y6_SIG_SIG ));
defparam clken_ctrl_X58_Y6_N1.coord_x = 14;
defparam clken_ctrl_X58_Y6_N1.coord_y = 9;
defparam clken_ctrl_X58_Y6_N1.coord_z = 1;
defparam clken_ctrl_X58_Y6_N1.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y6_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y7_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~62_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X58_Y7_SIG_SIG ));
defparam clken_ctrl_X58_Y7_N0.coord_x = 14;
defparam clken_ctrl_X58_Y7_N0.coord_y = 4;
defparam clken_ctrl_X58_Y7_N0.coord_z = 0;
defparam clken_ctrl_X58_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y7_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y7_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y7_SIG_VCC ));
defparam clken_ctrl_X58_Y7_N1.coord_x = 14;
defparam clken_ctrl_X58_Y7_N1.coord_y = 4;
defparam clken_ctrl_X58_Y7_N1.coord_z = 1;
defparam clken_ctrl_X58_Y7_N1.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y7_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X58_Y8_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~23_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y8_SIG_SIG ));
defparam clken_ctrl_X58_Y8_N0.coord_x = 17;
defparam clken_ctrl_X58_Y8_N0.coord_y = 5;
defparam clken_ctrl_X58_Y8_N0.coord_z = 0;
defparam clken_ctrl_X58_Y8_N0.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y8_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y8_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~65_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X58_Y8_SIG_SIG ));
defparam clken_ctrl_X58_Y8_N1.coord_x = 17;
defparam clken_ctrl_X58_Y8_N1.coord_y = 5;
defparam clken_ctrl_X58_Y8_N1.coord_z = 1;
defparam clken_ctrl_X58_Y8_N1.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y8_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y9_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~23_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y9_SIG_SIG ));
defparam clken_ctrl_X58_Y9_N0.coord_x = 18;
defparam clken_ctrl_X58_Y9_N0.coord_y = 9;
defparam clken_ctrl_X58_Y9_N0.coord_z = 0;
defparam clken_ctrl_X58_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y9_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X58_Y9_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~56_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X58_Y9_SIG_SIG ));
defparam clken_ctrl_X58_Y9_N1.coord_x = 18;
defparam clken_ctrl_X58_Y9_N1.coord_y = 9;
defparam clken_ctrl_X58_Y9_N1.coord_z = 1;
defparam clken_ctrl_X58_Y9_N1.ClkMux = 2'b10;
defparam clken_ctrl_X58_Y9_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y10_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~38_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X59_Y10_SIG_SIG ));
defparam clken_ctrl_X59_Y10_N0.coord_x = 18;
defparam clken_ctrl_X59_Y10_N0.coord_y = 6;
defparam clken_ctrl_X59_Y10_N0.coord_z = 0;
defparam clken_ctrl_X59_Y10_N0.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y10_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y10_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y10_SIG_VCC ));
defparam clken_ctrl_X59_Y10_N1.coord_x = 18;
defparam clken_ctrl_X59_Y10_N1.coord_y = 6;
defparam clken_ctrl_X59_Y10_N1.coord_z = 1;
defparam clken_ctrl_X59_Y10_N1.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y10_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X59_Y11_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~43_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X59_Y11_SIG_SIG ));
defparam clken_ctrl_X59_Y11_N0.coord_x = 19;
defparam clken_ctrl_X59_Y11_N0.coord_y = 3;
defparam clken_ctrl_X59_Y11_N0.coord_z = 0;
defparam clken_ctrl_X59_Y11_N0.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y11_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y11_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~34_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X59_Y11_SIG_SIG ));
defparam clken_ctrl_X59_Y11_N1.coord_x = 19;
defparam clken_ctrl_X59_Y11_N1.coord_y = 3;
defparam clken_ctrl_X59_Y11_N1.coord_z = 1;
defparam clken_ctrl_X59_Y11_N1.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y11_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y12_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~28_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X59_Y12_SIG_SIG ));
defparam clken_ctrl_X59_Y12_N0.coord_x = 20;
defparam clken_ctrl_X59_Y12_N0.coord_y = 5;
defparam clken_ctrl_X59_Y12_N0.coord_z = 0;
defparam clken_ctrl_X59_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y12_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y12_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y12_SIG_VCC ));
defparam clken_ctrl_X59_Y12_N1.coord_x = 20;
defparam clken_ctrl_X59_Y12_N1.coord_y = 5;
defparam clken_ctrl_X59_Y12_N1.coord_z = 1;
defparam clken_ctrl_X59_Y12_N1.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y12_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X59_Y1_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~72_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X59_Y1_SIG_SIG ));
defparam clken_ctrl_X59_Y1_N0.coord_x = 16;
defparam clken_ctrl_X59_Y1_N0.coord_y = 3;
defparam clken_ctrl_X59_Y1_N0.coord_z = 0;
defparam clken_ctrl_X59_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y1_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y1_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y1_SIG_VCC ));
defparam clken_ctrl_X59_Y1_N1.coord_x = 16;
defparam clken_ctrl_X59_Y1_N1.coord_y = 3;
defparam clken_ctrl_X59_Y1_N1.coord_z = 1;
defparam clken_ctrl_X59_Y1_N1.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y1_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X59_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~78_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X59_Y2_SIG_SIG ));
defparam clken_ctrl_X59_Y2_N0.coord_x = 10;
defparam clken_ctrl_X59_Y2_N0.coord_y = 3;
defparam clken_ctrl_X59_Y2_N0.coord_z = 0;
defparam clken_ctrl_X59_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y2_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y2_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y2_SIG_VCC ));
defparam clken_ctrl_X59_Y2_N1.coord_x = 10;
defparam clken_ctrl_X59_Y2_N1.coord_y = 3;
defparam clken_ctrl_X59_Y2_N1.coord_z = 1;
defparam clken_ctrl_X59_Y2_N1.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y2_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X59_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|Equal2~0_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X59_Y3_SIG_SIG ));
defparam clken_ctrl_X59_Y3_N0.coord_x = 15;
defparam clken_ctrl_X59_Y3_N0.coord_y = 12;
defparam clken_ctrl_X59_Y3_N0.coord_z = 0;
defparam clken_ctrl_X59_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y3_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y3_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y3_SIG_VCC ));
defparam clken_ctrl_X59_Y3_N1.coord_x = 15;
defparam clken_ctrl_X59_Y3_N1.coord_y = 12;
defparam clken_ctrl_X59_Y3_N1.coord_z = 1;
defparam clken_ctrl_X59_Y3_N1.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y3_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X59_Y4_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~45_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y4_SIG_SIG ));
defparam clken_ctrl_X59_Y4_N0.coord_x = 17;
defparam clken_ctrl_X59_Y4_N0.coord_y = 11;
defparam clken_ctrl_X59_Y4_N0.coord_z = 0;
defparam clken_ctrl_X59_Y4_N0.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y4_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y4_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~14_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X59_Y4_SIG_SIG ));
defparam clken_ctrl_X59_Y4_N1.coord_x = 17;
defparam clken_ctrl_X59_Y4_N1.coord_y = 11;
defparam clken_ctrl_X59_Y4_N1.coord_z = 1;
defparam clken_ctrl_X59_Y4_N1.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y4_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y5_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y5_SIG_VCC ));
defparam clken_ctrl_X59_Y5_N0.coord_x = 14;
defparam clken_ctrl_X59_Y5_N0.coord_y = 8;
defparam clken_ctrl_X59_Y5_N0.coord_z = 0;
defparam clken_ctrl_X59_Y5_N0.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y5_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X59_Y5_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~69_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X59_Y5_SIG_SIG ));
defparam clken_ctrl_X59_Y5_N1.coord_x = 14;
defparam clken_ctrl_X59_Y5_N1.coord_y = 8;
defparam clken_ctrl_X59_Y5_N1.coord_z = 1;
defparam clken_ctrl_X59_Y5_N1.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y5_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y6_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~49_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X59_Y6_SIG_SIG ));
defparam clken_ctrl_X59_Y6_N0.coord_x = 18;
defparam clken_ctrl_X59_Y6_N0.coord_y = 11;
defparam clken_ctrl_X59_Y6_N0.coord_z = 0;
defparam clken_ctrl_X59_Y6_N0.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y6_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y6_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|pwmUpdateTrigger~q ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|pwmUpdateTrigger~q_X59_Y6_SIG_SIG ));
defparam clken_ctrl_X59_Y6_N1.coord_x = 18;
defparam clken_ctrl_X59_Y6_N1.coord_y = 11;
defparam clken_ctrl_X59_Y6_N1.coord_z = 1;
defparam clken_ctrl_X59_Y6_N1.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y6_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y7_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~61_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X59_Y7_SIG_SIG ));
defparam clken_ctrl_X59_Y7_N0.coord_x = 18;
defparam clken_ctrl_X59_Y7_N0.coord_y = 5;
defparam clken_ctrl_X59_Y7_N0.coord_z = 0;
defparam clken_ctrl_X59_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y7_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y7_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~11_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X59_Y7_SIG_SIG ));
defparam clken_ctrl_X59_Y7_N1.coord_x = 18;
defparam clken_ctrl_X59_Y7_N1.coord_y = 5;
defparam clken_ctrl_X59_Y7_N1.coord_z = 1;
defparam clken_ctrl_X59_Y7_N1.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y7_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y8_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X59_Y8_SIG_SIG ));
defparam clken_ctrl_X59_Y8_N0.coord_x = 14;
defparam clken_ctrl_X59_Y8_N0.coord_y = 6;
defparam clken_ctrl_X59_Y8_N0.coord_z = 0;
defparam clken_ctrl_X59_Y8_N0.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y8_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y8_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~45_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y8_SIG_SIG ));
defparam clken_ctrl_X59_Y8_N1.coord_x = 14;
defparam clken_ctrl_X59_Y8_N1.coord_y = 6;
defparam clken_ctrl_X59_Y8_N1.coord_z = 1;
defparam clken_ctrl_X59_Y8_N1.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y8_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y9_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~25_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X59_Y9_SIG_SIG ));
defparam clken_ctrl_X59_Y9_N0.coord_x = 18;
defparam clken_ctrl_X59_Y9_N0.coord_y = 10;
defparam clken_ctrl_X59_Y9_N0.coord_z = 0;
defparam clken_ctrl_X59_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y9_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X59_Y9_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~49_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X59_Y9_SIG_SIG ));
defparam clken_ctrl_X59_Y9_N1.coord_x = 18;
defparam clken_ctrl_X59_Y9_N1.coord_y = 10;
defparam clken_ctrl_X59_Y9_N1.coord_z = 1;
defparam clken_ctrl_X59_Y9_N1.ClkMux = 2'b10;
defparam clken_ctrl_X59_Y9_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y10_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~66_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X60_Y10_SIG_SIG ));
defparam clken_ctrl_X60_Y10_N0.coord_x = 20;
defparam clken_ctrl_X60_Y10_N0.coord_y = 11;
defparam clken_ctrl_X60_Y10_N0.coord_z = 0;
defparam clken_ctrl_X60_Y10_N0.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y10_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y10_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~57_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X60_Y10_SIG_SIG ));
defparam clken_ctrl_X60_Y10_N1.coord_x = 20;
defparam clken_ctrl_X60_Y10_N1.coord_y = 11;
defparam clken_ctrl_X60_Y10_N1.coord_z = 1;
defparam clken_ctrl_X60_Y10_N1.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y10_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y11_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~34_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X60_Y11_SIG_SIG ));
defparam clken_ctrl_X60_Y11_N0.coord_x = 19;
defparam clken_ctrl_X60_Y11_N0.coord_y = 4;
defparam clken_ctrl_X60_Y11_N0.coord_z = 0;
defparam clken_ctrl_X60_Y11_N0.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y11_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y11_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~73_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X60_Y11_SIG_SIG ));
defparam clken_ctrl_X60_Y11_N1.coord_x = 19;
defparam clken_ctrl_X60_Y11_N1.coord_y = 4;
defparam clken_ctrl_X60_Y11_N1.coord_z = 1;
defparam clken_ctrl_X60_Y11_N1.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y11_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y12_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~28_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X60_Y12_SIG_SIG ));
defparam clken_ctrl_X60_Y12_N0.coord_x = 20;
defparam clken_ctrl_X60_Y12_N0.coord_y = 7;
defparam clken_ctrl_X60_Y12_N0.coord_z = 0;
defparam clken_ctrl_X60_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y12_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y12_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~38_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X60_Y12_SIG_SIG ));
defparam clken_ctrl_X60_Y12_N1.coord_x = 20;
defparam clken_ctrl_X60_Y12_N1.coord_y = 7;
defparam clken_ctrl_X60_Y12_N1.coord_z = 1;
defparam clken_ctrl_X60_Y12_N1.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y12_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y1_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~40_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X60_Y1_SIG_SIG ));
defparam clken_ctrl_X60_Y1_N0.coord_x = 17;
defparam clken_ctrl_X60_Y1_N0.coord_y = 1;
defparam clken_ctrl_X60_Y1_N0.coord_z = 0;
defparam clken_ctrl_X60_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y1_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y1_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X60_Y1_SIG_VCC ));
defparam clken_ctrl_X60_Y1_N1.coord_x = 17;
defparam clken_ctrl_X60_Y1_N1.coord_y = 1;
defparam clken_ctrl_X60_Y1_N1.coord_z = 1;
defparam clken_ctrl_X60_Y1_N1.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y1_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X60_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~52_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X60_Y2_SIG_SIG ));
defparam clken_ctrl_X60_Y2_N0.coord_x = 11;
defparam clken_ctrl_X60_Y2_N0.coord_y = 4;
defparam clken_ctrl_X60_Y2_N0.coord_z = 0;
defparam clken_ctrl_X60_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y2_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y2_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~31_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X60_Y2_SIG_SIG ));
defparam clken_ctrl_X60_Y2_N1.coord_x = 11;
defparam clken_ctrl_X60_Y2_N1.coord_y = 4;
defparam clken_ctrl_X60_Y2_N1.coord_z = 1;
defparam clken_ctrl_X60_Y2_N1.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y2_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|Equal2~0_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X60_Y3_SIG_SIG ));
defparam clken_ctrl_X60_Y3_N0.coord_x = 15;
defparam clken_ctrl_X60_Y3_N0.coord_y = 7;
defparam clken_ctrl_X60_Y3_N0.coord_z = 0;
defparam clken_ctrl_X60_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y3_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y3_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~80_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X60_Y3_SIG_SIG ));
defparam clken_ctrl_X60_Y3_N1.coord_x = 15;
defparam clken_ctrl_X60_Y3_N1.coord_y = 7;
defparam clken_ctrl_X60_Y3_N1.coord_z = 1;
defparam clken_ctrl_X60_Y3_N1.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y3_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y4_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~69_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X60_Y4_SIG_SIG ));
defparam clken_ctrl_X60_Y4_N0.coord_x = 15;
defparam clken_ctrl_X60_Y4_N0.coord_y = 8;
defparam clken_ctrl_X60_Y4_N0.coord_z = 0;
defparam clken_ctrl_X60_Y4_N0.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y4_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y4_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~11_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X60_Y4_SIG_SIG ));
defparam clken_ctrl_X60_Y4_N1.coord_x = 15;
defparam clken_ctrl_X60_Y4_N1.coord_y = 8;
defparam clken_ctrl_X60_Y4_N1.coord_z = 1;
defparam clken_ctrl_X60_Y4_N1.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y4_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y5_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~24_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X60_Y5_SIG_SIG ));
defparam clken_ctrl_X60_Y5_N0.coord_x = 15;
defparam clken_ctrl_X60_Y5_N0.coord_y = 10;
defparam clken_ctrl_X60_Y5_N0.coord_z = 0;
defparam clken_ctrl_X60_Y5_N0.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y5_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y5_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~59_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X60_Y5_SIG_SIG ));
defparam clken_ctrl_X60_Y5_N1.coord_x = 15;
defparam clken_ctrl_X60_Y5_N1.coord_y = 10;
defparam clken_ctrl_X60_Y5_N1.coord_z = 1;
defparam clken_ctrl_X60_Y5_N1.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y5_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y6_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~36_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X60_Y6_SIG_SIG ));
defparam clken_ctrl_X60_Y6_N0.coord_x = 18;
defparam clken_ctrl_X60_Y6_N0.coord_y = 7;
defparam clken_ctrl_X60_Y6_N0.coord_z = 0;
defparam clken_ctrl_X60_Y6_N0.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y6_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y6_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X60_Y6_SIG_VCC ));
defparam clken_ctrl_X60_Y6_N1.coord_x = 18;
defparam clken_ctrl_X60_Y6_N1.coord_y = 7;
defparam clken_ctrl_X60_Y6_N1.coord_z = 1;
defparam clken_ctrl_X60_Y6_N1.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y6_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X60_Y7_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~46_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X60_Y7_SIG_SIG ));
defparam clken_ctrl_X60_Y7_N0.coord_x = 18;
defparam clken_ctrl_X60_Y7_N0.coord_y = 4;
defparam clken_ctrl_X60_Y7_N0.coord_z = 0;
defparam clken_ctrl_X60_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y7_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y7_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~49_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X60_Y7_SIG_SIG ));
defparam clken_ctrl_X60_Y7_N1.coord_x = 18;
defparam clken_ctrl_X60_Y7_N1.coord_y = 4;
defparam clken_ctrl_X60_Y7_N1.coord_z = 1;
defparam clken_ctrl_X60_Y7_N1.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y7_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y8_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~42_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X60_Y8_SIG_SIG ));
defparam clken_ctrl_X60_Y8_N0.coord_x = 16;
defparam clken_ctrl_X60_Y8_N0.coord_y = 7;
defparam clken_ctrl_X60_Y8_N0.coord_z = 0;
defparam clken_ctrl_X60_Y8_N0.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y8_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y8_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~47_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X60_Y8_SIG_SIG ));
defparam clken_ctrl_X60_Y8_N1.coord_x = 16;
defparam clken_ctrl_X60_Y8_N1.coord_y = 7;
defparam clken_ctrl_X60_Y8_N1.coord_z = 1;
defparam clken_ctrl_X60_Y8_N1.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y8_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y9_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~43_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X60_Y9_SIG_SIG ));
defparam clken_ctrl_X60_Y9_N0.coord_x = 20;
defparam clken_ctrl_X60_Y9_N0.coord_y = 4;
defparam clken_ctrl_X60_Y9_N0.coord_z = 0;
defparam clken_ctrl_X60_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y9_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X60_Y9_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~60_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X60_Y9_SIG_SIG ));
defparam clken_ctrl_X60_Y9_N1.coord_x = 20;
defparam clken_ctrl_X60_Y9_N1.coord_y = 4;
defparam clken_ctrl_X60_Y9_N1.coord_z = 1;
defparam clken_ctrl_X60_Y9_N1.ClkMux = 2'b10;
defparam clken_ctrl_X60_Y9_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y10_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~36_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X61_Y10_SIG_SIG ));
defparam clken_ctrl_X61_Y10_N0.coord_x = 19;
defparam clken_ctrl_X61_Y10_N0.coord_y = 9;
defparam clken_ctrl_X61_Y10_N0.coord_z = 0;
defparam clken_ctrl_X61_Y10_N0.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y10_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y10_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~74_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X61_Y10_SIG_SIG ));
defparam clken_ctrl_X61_Y10_N1.coord_x = 19;
defparam clken_ctrl_X61_Y10_N1.coord_y = 9;
defparam clken_ctrl_X61_Y10_N1.coord_z = 1;
defparam clken_ctrl_X61_Y10_N1.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y10_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y11_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y11_SIG_VCC ));
defparam clken_ctrl_X61_Y11_N0.coord_x = 19;
defparam clken_ctrl_X61_Y11_N0.coord_y = 8;
defparam clken_ctrl_X61_Y11_N0.coord_z = 0;
defparam clken_ctrl_X61_Y11_N0.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y11_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X61_Y11_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~49_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X61_Y11_SIG_SIG ));
defparam clken_ctrl_X61_Y11_N1.coord_x = 19;
defparam clken_ctrl_X61_Y11_N1.coord_y = 8;
defparam clken_ctrl_X61_Y11_N1.coord_z = 1;
defparam clken_ctrl_X61_Y11_N1.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y11_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y12_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ));
defparam clken_ctrl_X61_Y12_N0.coord_x = 19;
defparam clken_ctrl_X61_Y12_N0.coord_y = 6;
defparam clken_ctrl_X61_Y12_N0.coord_z = 0;
defparam clken_ctrl_X61_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y12_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y12_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y12_SIG_VCC ));
defparam clken_ctrl_X61_Y12_N1.coord_x = 19;
defparam clken_ctrl_X61_Y12_N1.coord_y = 6;
defparam clken_ctrl_X61_Y12_N1.coord_z = 1;
defparam clken_ctrl_X61_Y12_N1.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y12_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X61_Y1_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y1_SIG_SIG ));
defparam clken_ctrl_X61_Y1_N0.coord_x = 18;
defparam clken_ctrl_X61_Y1_N0.coord_y = 1;
defparam clken_ctrl_X61_Y1_N0.coord_z = 0;
defparam clken_ctrl_X61_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y1_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y1_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~40_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X61_Y1_SIG_SIG ));
defparam clken_ctrl_X61_Y1_N1.coord_x = 18;
defparam clken_ctrl_X61_Y1_N1.coord_y = 1;
defparam clken_ctrl_X61_Y1_N1.coord_z = 1;
defparam clken_ctrl_X61_Y1_N1.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y1_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y2_SIG_VCC ));
defparam clken_ctrl_X61_Y2_N0.coord_x = 15;
defparam clken_ctrl_X61_Y2_N0.coord_y = 5;
defparam clken_ctrl_X61_Y2_N0.coord_z = 0;
defparam clken_ctrl_X61_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y2_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X61_Y2_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~80_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y2_SIG_SIG ));
defparam clken_ctrl_X61_Y2_N1.coord_x = 15;
defparam clken_ctrl_X61_Y2_N1.coord_y = 5;
defparam clken_ctrl_X61_Y2_N1.coord_z = 1;
defparam clken_ctrl_X61_Y2_N1.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y2_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~81_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X61_Y3_SIG_SIG ));
defparam clken_ctrl_X61_Y3_N0.coord_x = 15;
defparam clken_ctrl_X61_Y3_N0.coord_y = 1;
defparam clken_ctrl_X61_Y3_N0.coord_z = 0;
defparam clken_ctrl_X61_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y3_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y3_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~80_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y3_SIG_SIG ));
defparam clken_ctrl_X61_Y3_N1.coord_x = 15;
defparam clken_ctrl_X61_Y3_N1.coord_y = 1;
defparam clken_ctrl_X61_Y3_N1.coord_z = 1;
defparam clken_ctrl_X61_Y3_N1.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y3_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y4_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ));
defparam clken_ctrl_X61_Y4_N0.coord_x = 17;
defparam clken_ctrl_X61_Y4_N0.coord_y = 8;
defparam clken_ctrl_X61_Y4_N0.coord_z = 0;
defparam clken_ctrl_X61_Y4_N0.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y4_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X61_Y4_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~44_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X61_Y4_SIG_SIG ));
defparam clken_ctrl_X61_Y4_N1.coord_x = 17;
defparam clken_ctrl_X61_Y4_N1.coord_y = 8;
defparam clken_ctrl_X61_Y4_N1.coord_z = 1;
defparam clken_ctrl_X61_Y4_N1.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y4_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y5_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~31_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X61_Y5_SIG_SIG ));
defparam clken_ctrl_X61_Y5_N0.coord_x = 14;
defparam clken_ctrl_X61_Y5_N0.coord_y = 1;
defparam clken_ctrl_X61_Y5_N0.coord_z = 0;
defparam clken_ctrl_X61_Y5_N0.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y5_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y5_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y5_SIG_VCC ));
defparam clken_ctrl_X61_Y5_N1.coord_x = 14;
defparam clken_ctrl_X61_Y5_N1.coord_y = 1;
defparam clken_ctrl_X61_Y5_N1.coord_z = 1;
defparam clken_ctrl_X61_Y5_N1.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y5_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X61_Y6_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~64_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X61_Y6_SIG_SIG ));
defparam clken_ctrl_X61_Y6_N0.coord_x = 15;
defparam clken_ctrl_X61_Y6_N0.coord_y = 9;
defparam clken_ctrl_X61_Y6_N0.coord_z = 0;
defparam clken_ctrl_X61_Y6_N0.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y6_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y6_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~20_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X61_Y6_SIG_SIG ));
defparam clken_ctrl_X61_Y6_N1.coord_x = 15;
defparam clken_ctrl_X61_Y6_N1.coord_y = 9;
defparam clken_ctrl_X61_Y6_N1.coord_z = 1;
defparam clken_ctrl_X61_Y6_N1.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y6_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y7_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~46_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X61_Y7_SIG_SIG ));
defparam clken_ctrl_X61_Y7_N0.coord_x = 17;
defparam clken_ctrl_X61_Y7_N0.coord_y = 3;
defparam clken_ctrl_X61_Y7_N0.coord_z = 0;
defparam clken_ctrl_X61_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y7_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y7_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~77_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X61_Y7_SIG_SIG ));
defparam clken_ctrl_X61_Y7_N1.coord_x = 17;
defparam clken_ctrl_X61_Y7_N1.coord_y = 3;
defparam clken_ctrl_X61_Y7_N1.coord_z = 1;
defparam clken_ctrl_X61_Y7_N1.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y7_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y8_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~73_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X61_Y8_SIG_SIG ));
defparam clken_ctrl_X61_Y8_N0.coord_x = 19;
defparam clken_ctrl_X61_Y8_N0.coord_y = 2;
defparam clken_ctrl_X61_Y8_N0.coord_z = 0;
defparam clken_ctrl_X61_Y8_N0.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y8_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X61_Y8_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y8_SIG_VCC ));
defparam clken_ctrl_X61_Y8_N1.coord_x = 19;
defparam clken_ctrl_X61_Y8_N1.coord_y = 2;
defparam clken_ctrl_X61_Y8_N1.coord_z = 1;
defparam clken_ctrl_X61_Y8_N1.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y8_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X61_Y9_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y9_SIG_VCC ));
defparam clken_ctrl_X61_Y9_N0.coord_x = 19;
defparam clken_ctrl_X61_Y9_N0.coord_y = 7;
defparam clken_ctrl_X61_Y9_N0.coord_z = 0;
defparam clken_ctrl_X61_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y9_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X61_Y9_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~60_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X61_Y9_SIG_SIG ));
defparam clken_ctrl_X61_Y9_N1.coord_x = 19;
defparam clken_ctrl_X61_Y9_N1.coord_y = 7;
defparam clken_ctrl_X61_Y9_N1.coord_z = 1;
defparam clken_ctrl_X61_Y9_N1.ClkMux = 2'b10;
defparam clken_ctrl_X61_Y9_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y10_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y10_SIG_VCC ));
defparam clken_ctrl_X62_Y10_N0.coord_x = 20;
defparam clken_ctrl_X62_Y10_N0.coord_y = 12;
defparam clken_ctrl_X62_Y10_N0.coord_z = 0;
defparam clken_ctrl_X62_Y10_N0.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y10_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X62_Y10_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~74_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X62_Y10_SIG_SIG ));
defparam clken_ctrl_X62_Y10_N1.coord_x = 20;
defparam clken_ctrl_X62_Y10_N1.coord_y = 12;
defparam clken_ctrl_X62_Y10_N1.coord_z = 1;
defparam clken_ctrl_X62_Y10_N1.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y10_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y11_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y11_SIG_SIG ));
defparam clken_ctrl_X62_Y11_N0.coord_x = 20;
defparam clken_ctrl_X62_Y11_N0.coord_y = 9;
defparam clken_ctrl_X62_Y11_N0.coord_z = 0;
defparam clken_ctrl_X62_Y11_N0.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y11_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y11_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~68_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y11_SIG_SIG ));
defparam clken_ctrl_X62_Y11_N1.coord_x = 20;
defparam clken_ctrl_X62_Y11_N1.coord_y = 9;
defparam clken_ctrl_X62_Y11_N1.coord_z = 1;
defparam clken_ctrl_X62_Y11_N1.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y11_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y12_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ));
defparam clken_ctrl_X62_Y12_N0.coord_x = 20;
defparam clken_ctrl_X62_Y12_N0.coord_y = 6;
defparam clken_ctrl_X62_Y12_N0.coord_z = 0;
defparam clken_ctrl_X62_Y12_N0.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y12_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y12_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y12_SIG_VCC ));
defparam clken_ctrl_X62_Y12_N1.coord_x = 20;
defparam clken_ctrl_X62_Y12_N1.coord_y = 6;
defparam clken_ctrl_X62_Y12_N1.coord_z = 1;
defparam clken_ctrl_X62_Y12_N1.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y12_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X62_Y1_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~81_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X62_Y1_SIG_SIG ));
defparam clken_ctrl_X62_Y1_N0.coord_x = 12;
defparam clken_ctrl_X62_Y1_N0.coord_y = 1;
defparam clken_ctrl_X62_Y1_N0.coord_z = 0;
defparam clken_ctrl_X62_Y1_N0.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y1_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y1_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y1_SIG_VCC ));
defparam clken_ctrl_X62_Y1_N1.coord_x = 12;
defparam clken_ctrl_X62_Y1_N1.coord_y = 1;
defparam clken_ctrl_X62_Y1_N1.coord_z = 1;
defparam clken_ctrl_X62_Y1_N1.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y1_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X62_Y2_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y2_SIG_SIG ));
defparam clken_ctrl_X62_Y2_N0.coord_x = 17;
defparam clken_ctrl_X62_Y2_N0.coord_y = 6;
defparam clken_ctrl_X62_Y2_N0.coord_z = 0;
defparam clken_ctrl_X62_Y2_N0.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y2_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y2_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~44_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X62_Y2_SIG_SIG ));
defparam clken_ctrl_X62_Y2_N1.coord_x = 17;
defparam clken_ctrl_X62_Y2_N1.coord_y = 6;
defparam clken_ctrl_X62_Y2_N1.coord_z = 1;
defparam clken_ctrl_X62_Y2_N1.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y2_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y3_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y3_SIG_VCC ));
defparam clken_ctrl_X62_Y3_N0.coord_x = 16;
defparam clken_ctrl_X62_Y3_N0.coord_y = 6;
defparam clken_ctrl_X62_Y3_N0.coord_z = 0;
defparam clken_ctrl_X62_Y3_N0.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y3_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X62_Y3_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~77_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X62_Y3_SIG_SIG ));
defparam clken_ctrl_X62_Y3_N1.coord_x = 16;
defparam clken_ctrl_X62_Y3_N1.coord_y = 6;
defparam clken_ctrl_X62_Y3_N1.coord_z = 1;
defparam clken_ctrl_X62_Y3_N1.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y3_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y4_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~47_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X62_Y4_SIG_SIG ));
defparam clken_ctrl_X62_Y4_N0.coord_x = 14;
defparam clken_ctrl_X62_Y4_N0.coord_y = 3;
defparam clken_ctrl_X62_Y4_N0.coord_z = 0;
defparam clken_ctrl_X62_Y4_N0.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y4_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y4_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y4_SIG_VCC ));
defparam clken_ctrl_X62_Y4_N1.coord_x = 14;
defparam clken_ctrl_X62_Y4_N1.coord_y = 3;
defparam clken_ctrl_X62_Y4_N1.coord_z = 1;
defparam clken_ctrl_X62_Y4_N1.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y4_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X62_Y5_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y5_SIG_VCC ));
defparam clken_ctrl_X62_Y5_N0.coord_x = 17;
defparam clken_ctrl_X62_Y5_N0.coord_y = 10;
defparam clken_ctrl_X62_Y5_N0.coord_z = 0;
defparam clken_ctrl_X62_Y5_N0.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y5_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X62_Y5_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~64_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X62_Y5_SIG_SIG ));
defparam clken_ctrl_X62_Y5_N1.coord_x = 17;
defparam clken_ctrl_X62_Y5_N1.coord_y = 10;
defparam clken_ctrl_X62_Y5_N1.coord_z = 1;
defparam clken_ctrl_X62_Y5_N1.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y5_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y6_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~20_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X62_Y6_SIG_SIG ));
defparam clken_ctrl_X62_Y6_N0.coord_x = 17;
defparam clken_ctrl_X62_Y6_N0.coord_y = 12;
defparam clken_ctrl_X62_Y6_N0.coord_z = 0;
defparam clken_ctrl_X62_Y6_N0.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y6_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y6_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~42_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X62_Y6_SIG_SIG ));
defparam clken_ctrl_X62_Y6_N1.coord_x = 17;
defparam clken_ctrl_X62_Y6_N1.coord_y = 12;
defparam clken_ctrl_X62_Y6_N1.coord_z = 1;
defparam clken_ctrl_X62_Y6_N1.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y6_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y7_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y7_SIG_VCC ));
defparam clken_ctrl_X62_Y7_N0.coord_x = 15;
defparam clken_ctrl_X62_Y7_N0.coord_y = 6;
defparam clken_ctrl_X62_Y7_N0.coord_z = 0;
defparam clken_ctrl_X62_Y7_N0.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y7_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X62_Y7_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~68_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y7_SIG_SIG ));
defparam clken_ctrl_X62_Y7_N1.coord_x = 15;
defparam clken_ctrl_X62_Y7_N1.coord_y = 6;
defparam clken_ctrl_X62_Y7_N1.coord_z = 1;
defparam clken_ctrl_X62_Y7_N1.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y7_N1.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y8_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~33_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X62_Y8_SIG_SIG ));
defparam clken_ctrl_X62_Y8_N0.coord_x = 18;
defparam clken_ctrl_X62_Y8_N0.coord_y = 2;
defparam clken_ctrl_X62_Y8_N0.coord_z = 0;
defparam clken_ctrl_X62_Y8_N0.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y8_N0.ClkEnMux = 2'b10;

alta_clkenctrl clken_ctrl_X62_Y8_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y8_SIG_VCC ));
defparam clken_ctrl_X62_Y8_N1.coord_x = 18;
defparam clken_ctrl_X62_Y8_N1.coord_y = 2;
defparam clken_ctrl_X62_Y8_N1.coord_z = 1;
defparam clken_ctrl_X62_Y8_N1.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y8_N1.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X62_Y9_N0(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y9_SIG_VCC ));
defparam clken_ctrl_X62_Y9_N0.coord_x = 19;
defparam clken_ctrl_X62_Y9_N0.coord_y = 11;
defparam clken_ctrl_X62_Y9_N0.coord_z = 0;
defparam clken_ctrl_X62_Y9_N0.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y9_N0.ClkEnMux = 2'b01;

alta_clkenctrl clken_ctrl_X62_Y9_N1(
	.ClkIn(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ),
	.ClkEn(\macro_inst|controller|sm_pwm|Decoder0~66_combout ),
	.ClkOut(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X62_Y9_SIG_SIG ));
defparam clken_ctrl_X62_Y9_N1.coord_x = 19;
defparam clken_ctrl_X62_Y9_N1.coord_y = 11;
defparam clken_ctrl_X62_Y9_N1.coord_z = 1;
defparam clken_ctrl_X62_Y9_N1.ClkMux = 2'b10;
defparam clken_ctrl_X62_Y9_N1.ClkEnMux = 2'b10;

alta_io_gclk \gclksw_inst|gclk_switch (
	.inclk(\gclksw_inst|gclk_switch__alta_gclksw__clkout ),
	.outclk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp ));
defparam \gclksw_inst|gclk_switch .coord_x = 22;
defparam \gclksw_inst|gclk_switch .coord_y = 4;
defparam \gclksw_inst|gclk_switch .coord_z = 5;

alta_gclksw \gclksw_inst|gclk_switch__alta_gclksw (
	.resetn(\rv32.resetn_out ),
	.clkin0(\PIN_HSI~input_o ),
	.clkin1(\PIN_HSE~input_o ),
	.clkin2(\pll_inst|auto_generated|pll1_CLK_bus [0]),
	.clkin3(1'bx),
	.select({\rv32.sys_ctrl_clkSource[1] , \rv32.sys_ctrl_clkSource[0] }),
	.clkout(\gclksw_inst|gclk_switch__alta_gclksw__clkout ));
defparam \gclksw_inst|gclk_switch__alta_gclksw .coord_x = 22;
defparam \gclksw_inst|gclk_switch__alta_gclksw .coord_y = 4;
defparam \gclksw_inst|gclk_switch__alta_gclksw .coord_z = 0;

alta_slice \macro_inst|Add0~10 (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~10_combout ),
	.Cout(\macro_inst|Add0~11 ),
	.Q());
defparam \macro_inst|Add0~10 .coord_x = 3;
defparam \macro_inst|Add0~10 .coord_y = 2;
defparam \macro_inst|Add0~10 .coord_z = 10;
defparam \macro_inst|Add0~10 .mask = 16'h3C3F;
defparam \macro_inst|Add0~10 .modeMux = 1'b1;
defparam \macro_inst|Add0~10 .FeedbackMux = 1'b0;
defparam \macro_inst|Add0~10 .ShiftMux = 1'b0;
defparam \macro_inst|Add0~10 .BypassEn = 1'b0;
defparam \macro_inst|Add0~10 .CarryEnb = 1'b0;

alta_slice \macro_inst|Add0~14 (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~14_combout ),
	.Cout(\macro_inst|Add0~15 ),
	.Q());
defparam \macro_inst|Add0~14 .coord_x = 3;
defparam \macro_inst|Add0~14 .coord_y = 2;
defparam \macro_inst|Add0~14 .coord_z = 12;
defparam \macro_inst|Add0~14 .mask = 16'h3C3F;
defparam \macro_inst|Add0~14 .modeMux = 1'b1;
defparam \macro_inst|Add0~14 .FeedbackMux = 1'b0;
defparam \macro_inst|Add0~14 .ShiftMux = 1'b0;
defparam \macro_inst|Add0~14 .BypassEn = 1'b0;
defparam \macro_inst|Add0~14 .CarryEnb = 1'b0;

alta_slice \macro_inst|Add0~16 (
	.A(\macro_inst|clk10hz_cnt [8]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~15 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~16_combout ),
	.Cout(\macro_inst|Add0~17 ),
	.Q());
defparam \macro_inst|Add0~16 .coord_x = 3;
defparam \macro_inst|Add0~16 .coord_y = 2;
defparam \macro_inst|Add0~16 .coord_z = 13;
defparam \macro_inst|Add0~16 .mask = 16'hA50A;
defparam \macro_inst|Add0~16 .modeMux = 1'b1;
defparam \macro_inst|Add0~16 .FeedbackMux = 1'b0;
defparam \macro_inst|Add0~16 .ShiftMux = 1'b0;
defparam \macro_inst|Add0~16 .BypassEn = 1'b0;
defparam \macro_inst|Add0~16 .CarryEnb = 1'b0;

alta_slice \macro_inst|Add0~18 (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [9]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~17 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~18_combout ),
	.Cout(\macro_inst|Add0~19 ),
	.Q());
defparam \macro_inst|Add0~18 .coord_x = 3;
defparam \macro_inst|Add0~18 .coord_y = 2;
defparam \macro_inst|Add0~18 .coord_z = 14;
defparam \macro_inst|Add0~18 .mask = 16'h3C3F;
defparam \macro_inst|Add0~18 .modeMux = 1'b1;
defparam \macro_inst|Add0~18 .FeedbackMux = 1'b0;
defparam \macro_inst|Add0~18 .ShiftMux = 1'b0;
defparam \macro_inst|Add0~18 .BypassEn = 1'b0;
defparam \macro_inst|Add0~18 .CarryEnb = 1'b0;

alta_slice \macro_inst|Add0~20 (
	.A(\macro_inst|clk10hz_cnt [10]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~19 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~20_combout ),
	.Cout(\macro_inst|Add0~21 ),
	.Q());
defparam \macro_inst|Add0~20 .coord_x = 3;
defparam \macro_inst|Add0~20 .coord_y = 2;
defparam \macro_inst|Add0~20 .coord_z = 15;
defparam \macro_inst|Add0~20 .mask = 16'hA50A;
defparam \macro_inst|Add0~20 .modeMux = 1'b1;
defparam \macro_inst|Add0~20 .FeedbackMux = 1'b0;
defparam \macro_inst|Add0~20 .ShiftMux = 1'b0;
defparam \macro_inst|Add0~20 .BypassEn = 1'b0;
defparam \macro_inst|Add0~20 .CarryEnb = 1'b0;

alta_slice \macro_inst|Add0~22 (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [11]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~21 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~22_combout ),
	.Cout(\macro_inst|Add0~23 ),
	.Q());
defparam \macro_inst|Add0~22 .coord_x = 3;
defparam \macro_inst|Add0~22 .coord_y = 1;
defparam \macro_inst|Add0~22 .coord_z = 0;
defparam \macro_inst|Add0~22 .mask = 16'h3C3F;
defparam \macro_inst|Add0~22 .modeMux = 1'b1;
defparam \macro_inst|Add0~22 .FeedbackMux = 1'b0;
defparam \macro_inst|Add0~22 .ShiftMux = 1'b0;
defparam \macro_inst|Add0~22 .BypassEn = 1'b0;
defparam \macro_inst|Add0~22 .CarryEnb = 1'b0;

alta_slice \macro_inst|Equal1~0 (
	.A(\rv32.mem_ahb_haddr[5] ),
	.B(\rv32.mem_ahb_haddr[12] ),
	.C(\rv32.mem_ahb_haddr[30] ),
	.D(\rv32.mem_ahb_haddr[29] ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal1~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal1~0 .coord_x = 14;
defparam \macro_inst|Equal1~0 .coord_y = 11;
defparam \macro_inst|Equal1~0 .coord_z = 2;
defparam \macro_inst|Equal1~0 .mask = 16'h4000;
defparam \macro_inst|Equal1~0 .modeMux = 1'b0;
defparam \macro_inst|Equal1~0 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal1~0 .ShiftMux = 1'b0;
defparam \macro_inst|Equal1~0 .BypassEn = 1'b0;
defparam \macro_inst|Equal1~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal1~1 (
	.A(\rv32.mem_ahb_haddr[23] ),
	.B(\rv32.mem_ahb_haddr[21] ),
	.C(\rv32.mem_ahb_haddr[9] ),
	.D(\rv32.mem_ahb_haddr[10] ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal1~1_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal1~1 .coord_x = 16;
defparam \macro_inst|Equal1~1 .coord_y = 11;
defparam \macro_inst|Equal1~1 .coord_z = 7;
defparam \macro_inst|Equal1~1 .mask = 16'h0001;
defparam \macro_inst|Equal1~1 .modeMux = 1'b0;
defparam \macro_inst|Equal1~1 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal1~1 .ShiftMux = 1'b0;
defparam \macro_inst|Equal1~1 .BypassEn = 1'b0;
defparam \macro_inst|Equal1~1 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal1~2 (
	.A(\rv32.mem_ahb_haddr[13] ),
	.B(\rv32.mem_ahb_haddr[28] ),
	.C(\rv32.mem_ahb_haddr[19] ),
	.D(\rv32.mem_ahb_haddr[8] ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal1~2_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal1~2 .coord_x = 14;
defparam \macro_inst|Equal1~2 .coord_y = 11;
defparam \macro_inst|Equal1~2 .coord_z = 6;
defparam \macro_inst|Equal1~2 .mask = 16'h0001;
defparam \macro_inst|Equal1~2 .modeMux = 1'b0;
defparam \macro_inst|Equal1~2 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal1~2 .ShiftMux = 1'b0;
defparam \macro_inst|Equal1~2 .BypassEn = 1'b0;
defparam \macro_inst|Equal1~2 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal1~3 (
	.A(\rv32.mem_ahb_haddr[25] ),
	.B(\rv32.mem_ahb_haddr[26] ),
	.C(\rv32.mem_ahb_haddr[20] ),
	.D(\rv32.mem_ahb_haddr[14] ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal1~3_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal1~3 .coord_x = 14;
defparam \macro_inst|Equal1~3 .coord_y = 11;
defparam \macro_inst|Equal1~3 .coord_z = 9;
defparam \macro_inst|Equal1~3 .mask = 16'h0001;
defparam \macro_inst|Equal1~3 .modeMux = 1'b0;
defparam \macro_inst|Equal1~3 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal1~3 .ShiftMux = 1'b0;
defparam \macro_inst|Equal1~3 .BypassEn = 1'b0;
defparam \macro_inst|Equal1~3 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal1~4 (
	.A(\macro_inst|Equal1~0_combout ),
	.B(\macro_inst|Equal1~3_combout ),
	.C(\macro_inst|Equal1~2_combout ),
	.D(\macro_inst|Equal1~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal1~4_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal1~4 .coord_x = 14;
defparam \macro_inst|Equal1~4 .coord_y = 11;
defparam \macro_inst|Equal1~4 .coord_z = 12;
defparam \macro_inst|Equal1~4 .mask = 16'h8000;
defparam \macro_inst|Equal1~4 .modeMux = 1'b0;
defparam \macro_inst|Equal1~4 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal1~4 .ShiftMux = 1'b0;
defparam \macro_inst|Equal1~4 .BypassEn = 1'b0;
defparam \macro_inst|Equal1~4 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal1~6 (
	.A(\rv32.mem_ahb_haddr[16] ),
	.B(\rv32.mem_ahb_haddr[7] ),
	.C(\rv32.mem_ahb_haddr[15] ),
	.D(\rv32.mem_ahb_haddr[6] ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal1~6_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal1~6 .coord_x = 15;
defparam \macro_inst|Equal1~6 .coord_y = 11;
defparam \macro_inst|Equal1~6 .coord_z = 14;
defparam \macro_inst|Equal1~6 .mask = 16'h0001;
defparam \macro_inst|Equal1~6 .modeMux = 1'b0;
defparam \macro_inst|Equal1~6 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal1~6 .ShiftMux = 1'b0;
defparam \macro_inst|Equal1~6 .BypassEn = 1'b0;
defparam \macro_inst|Equal1~6 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal1~7 (
	.A(\rv32.mem_ahb_haddr[4] ),
	.B(\rv32.mem_ahb_haddr[24] ),
	.C(\rv32.mem_ahb_haddr[22] ),
	.D(\rv32.mem_ahb_haddr[11] ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal1~7_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal1~7 .coord_x = 14;
defparam \macro_inst|Equal1~7 .coord_y = 11;
defparam \macro_inst|Equal1~7 .coord_z = 0;
defparam \macro_inst|Equal1~7 .mask = 16'h0001;
defparam \macro_inst|Equal1~7 .modeMux = 1'b0;
defparam \macro_inst|Equal1~7 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal1~7 .ShiftMux = 1'b0;
defparam \macro_inst|Equal1~7 .BypassEn = 1'b0;
defparam \macro_inst|Equal1~7 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal1~8 (
	.A(\macro_inst|Equal1~5_combout ),
	.B(\macro_inst|Equal1~6_combout ),
	.C(\macro_inst|Equal1~7_combout ),
	.D(\macro_inst|Equal1~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal1~8_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal1~8 .coord_x = 15;
defparam \macro_inst|Equal1~8 .coord_y = 11;
defparam \macro_inst|Equal1~8 .coord_z = 15;
defparam \macro_inst|Equal1~8 .mask = 16'h8000;
defparam \macro_inst|Equal1~8 .modeMux = 1'b0;
defparam \macro_inst|Equal1~8 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal1~8 .ShiftMux = 1'b0;
defparam \macro_inst|Equal1~8 .BypassEn = 1'b0;
defparam \macro_inst|Equal1~8 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal2~0 (
	.A(vcc),
	.B(vcc),
	.C(\rv32.mem_ahb_htrans[1] ),
	.D(\rv32.mem_ahb_htrans[0] ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal2~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal2~0 .coord_x = 14;
defparam \macro_inst|Equal2~0 .coord_y = 11;
defparam \macro_inst|Equal2~0 .coord_z = 14;
defparam \macro_inst|Equal2~0 .mask = 16'h00F0;
defparam \macro_inst|Equal2~0 .modeMux = 1'b0;
defparam \macro_inst|Equal2~0 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal2~0 .ShiftMux = 1'b0;
defparam \macro_inst|Equal2~0 .BypassEn = 1'b0;
defparam \macro_inst|Equal2~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal3~0 (
	.A(\macro_inst|clk10hz_cnt [19]),
	.B(\macro_inst|clk10hz_cnt [20]),
	.C(\macro_inst|clk10hz_cnt [21]),
	.D(\macro_inst|clk10hz_cnt [22]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal3~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal3~0 .coord_x = 3;
defparam \macro_inst|Equal3~0 .coord_y = 1;
defparam \macro_inst|Equal3~0 .coord_z = 14;
defparam \macro_inst|Equal3~0 .mask = 16'h0001;
defparam \macro_inst|Equal3~0 .modeMux = 1'b0;
defparam \macro_inst|Equal3~0 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal3~0 .ShiftMux = 1'b0;
defparam \macro_inst|Equal3~0 .BypassEn = 1'b0;
defparam \macro_inst|Equal3~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal3~1 (
	.A(\macro_inst|clk10hz_cnt [17]),
	.B(\macro_inst|clk10hz_cnt [18]),
	.C(\macro_inst|clk10hz_cnt [15]),
	.D(\macro_inst|clk10hz_cnt [16]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal3~1_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal3~1 .coord_x = 3;
defparam \macro_inst|Equal3~1 .coord_y = 1;
defparam \macro_inst|Equal3~1 .coord_z = 12;
defparam \macro_inst|Equal3~1 .mask = 16'h0001;
defparam \macro_inst|Equal3~1 .modeMux = 1'b0;
defparam \macro_inst|Equal3~1 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal3~1 .ShiftMux = 1'b0;
defparam \macro_inst|Equal3~1 .BypassEn = 1'b0;
defparam \macro_inst|Equal3~1 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal3~2 (
	.A(\macro_inst|clk10hz_cnt [11]),
	.B(\macro_inst|clk10hz_cnt [12]),
	.C(\macro_inst|clk10hz_cnt [13]),
	.D(\macro_inst|clk10hz_cnt [14]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal3~2_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal3~2 .coord_x = 3;
defparam \macro_inst|Equal3~2 .coord_y = 1;
defparam \macro_inst|Equal3~2 .coord_z = 13;
defparam \macro_inst|Equal3~2 .mask = 16'h0002;
defparam \macro_inst|Equal3~2 .modeMux = 1'b0;
defparam \macro_inst|Equal3~2 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal3~2 .ShiftMux = 1'b0;
defparam \macro_inst|Equal3~2 .BypassEn = 1'b0;
defparam \macro_inst|Equal3~2 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal3~3 (
	.A(\macro_inst|clk10hz_cnt [10]),
	.B(\macro_inst|clk10hz_cnt [9]),
	.C(\macro_inst|clk10hz_cnt [8]),
	.D(\macro_inst|clk10hz_cnt [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal3~3_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal3~3 .coord_x = 4;
defparam \macro_inst|Equal3~3 .coord_y = 2;
defparam \macro_inst|Equal3~3 .coord_z = 2;
defparam \macro_inst|Equal3~3 .mask = 16'h8000;
defparam \macro_inst|Equal3~3 .modeMux = 1'b0;
defparam \macro_inst|Equal3~3 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal3~3 .ShiftMux = 1'b0;
defparam \macro_inst|Equal3~3 .BypassEn = 1'b0;
defparam \macro_inst|Equal3~3 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal3~4 (
	.A(\macro_inst|Equal3~3_combout ),
	.B(\macro_inst|Equal3~1_combout ),
	.C(\macro_inst|Equal3~0_combout ),
	.D(\macro_inst|Equal3~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal3~4_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal3~4 .coord_x = 4;
defparam \macro_inst|Equal3~4 .coord_y = 2;
defparam \macro_inst|Equal3~4 .coord_z = 11;
defparam \macro_inst|Equal3~4 .mask = 16'h8000;
defparam \macro_inst|Equal3~4 .modeMux = 1'b0;
defparam \macro_inst|Equal3~4 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal3~4 .ShiftMux = 1'b0;
defparam \macro_inst|Equal3~4 .BypassEn = 1'b0;
defparam \macro_inst|Equal3~4 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal3~5 (
	.A(\macro_inst|clk10hz_cnt [5]),
	.B(\macro_inst|clk10hz_cnt [6]),
	.C(\macro_inst|clk10hz_cnt [3]),
	.D(\macro_inst|clk10hz_cnt [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal3~5_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal3~5 .coord_x = 3;
defparam \macro_inst|Equal3~5 .coord_y = 2;
defparam \macro_inst|Equal3~5 .coord_z = 2;
defparam \macro_inst|Equal3~5 .mask = 16'h1000;
defparam \macro_inst|Equal3~5 .modeMux = 1'b0;
defparam \macro_inst|Equal3~5 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal3~5 .ShiftMux = 1'b0;
defparam \macro_inst|Equal3~5 .BypassEn = 1'b0;
defparam \macro_inst|Equal3~5 .CarryEnb = 1'b1;

alta_slice \macro_inst|Equal3~6 (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [1]),
	.C(\macro_inst|clk10hz_cnt [0]),
	.D(\macro_inst|clk10hz_cnt [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Equal3~6_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|Equal3~6 .coord_x = 4;
defparam \macro_inst|Equal3~6 .coord_y = 4;
defparam \macro_inst|Equal3~6 .coord_z = 0;
defparam \macro_inst|Equal3~6 .mask = 16'hC000;
defparam \macro_inst|Equal3~6 .modeMux = 1'b0;
defparam \macro_inst|Equal3~6 .FeedbackMux = 1'b0;
defparam \macro_inst|Equal3~6 .ShiftMux = 1'b0;
defparam \macro_inst|Equal3~6 .BypassEn = 1'b0;
defparam \macro_inst|Equal3~6 .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[10] (
	.A(\macro_inst|ahb_add_reg [9]),
	.B(\macro_inst|ahb_add_reg [11]),
	.C(\rv32.mem_ahb_haddr[10] ),
	.D(\macro_inst|ahb_add_reg [8]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [10]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X59_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y3_SIG ),
	.SyncReset(SyncReset_X59_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Equal0~0_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [10]));
defparam \macro_inst|ahb_add_reg[10] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[10] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[10] .coord_z = 2;
defparam \macro_inst|ahb_add_reg[10] .mask = 16'h0100;
defparam \macro_inst|ahb_add_reg[10] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[10] .FeedbackMux = 1'b1;
defparam \macro_inst|ahb_add_reg[10] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[10] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[10] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[11] (
	.A(\macro_inst|ahb_add_reg [6]),
	.B(\macro_inst|ahb_add_reg [4]),
	.C(\rv32.mem_ahb_haddr[11] ),
	.D(\macro_inst|ahb_add_reg [5]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [11]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X59_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y3_SIG ),
	.SyncReset(SyncReset_X59_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~55_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [11]));
defparam \macro_inst|ahb_add_reg[11] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[11] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[11] .coord_z = 9;
defparam \macro_inst|ahb_add_reg[11] .mask = 16'h4400;
defparam \macro_inst|ahb_add_reg[11] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[11] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[11] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[11] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[11] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[12] (
	.A(\macro_inst|ahb_add_reg [15]),
	.B(\macro_inst|ahb_add_reg [13]),
	.C(\rv32.mem_ahb_haddr[12] ),
	.D(\macro_inst|ahb_add_reg [14]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [12]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X59_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y3_SIG ),
	.SyncReset(SyncReset_X59_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan0~0_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [12]));
defparam \macro_inst|ahb_add_reg[12] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[12] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[12] .coord_z = 8;
defparam \macro_inst|ahb_add_reg[12] .mask = 16'h0001;
defparam \macro_inst|ahb_add_reg[12] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[12] .FeedbackMux = 1'b1;
defparam \macro_inst|ahb_add_reg[12] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[12] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[12] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[13] (
	.A(\macro_inst|ahb_add_reg [6]),
	.B(\macro_inst|ahb_add_reg [4]),
	.C(\rv32.mem_ahb_haddr[13] ),
	.D(\macro_inst|ahb_add_reg [5]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [13]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X59_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y3_SIG ),
	.SyncReset(SyncReset_X59_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~51_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [13]));
defparam \macro_inst|ahb_add_reg[13] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[13] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[13] .coord_z = 3;
defparam \macro_inst|ahb_add_reg[13] .mask = 16'h1100;
defparam \macro_inst|ahb_add_reg[13] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[13] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[13] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[13] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[13] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[14] (
	.A(vcc),
	.B(\macro_inst|ahb_add_reg [7]),
	.C(\rv32.mem_ahb_haddr[14] ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~7_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [14]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X59_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y3_SIG ),
	.SyncReset(SyncReset_X59_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~8_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [14]));
defparam \macro_inst|ahb_add_reg[14] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[14] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[14] .coord_z = 4;
defparam \macro_inst|ahb_add_reg[14] .mask = 16'h3300;
defparam \macro_inst|ahb_add_reg[14] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[14] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[14] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[14] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[14] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[15] (
	.A(\macro_inst|ahb_add_reg [6]),
	.B(\macro_inst|ahb_add_reg [5]),
	.C(\rv32.mem_ahb_haddr[15] ),
	.D(\macro_inst|ahb_add_reg [7]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [15]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X59_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y3_SIG ),
	.SyncReset(SyncReset_X59_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Equal0~1_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [15]));
defparam \macro_inst|ahb_add_reg[15] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[15] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[15] .coord_z = 11;
defparam \macro_inst|ahb_add_reg[15] .mask = 16'h8800;
defparam \macro_inst|ahb_add_reg[15] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[15] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[15] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[15] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[15] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[16] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [16]),
	.C(\rv32.mem_ahb_haddr[16] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [16]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X58_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y3_SIG ),
	.SyncReset(SyncReset_X58_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y3_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[16]~16_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [16]));
defparam \macro_inst|ahb_add_reg[16] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[16] .coord_y = 11;
defparam \macro_inst|ahb_add_reg[16] .coord_z = 0;
defparam \macro_inst|ahb_add_reg[16] .mask = 16'hCC00;
defparam \macro_inst|ahb_add_reg[16] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[16] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[16] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[16] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[16] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[17] (
	.A(\macro_inst|ahb_add_reg [20]),
	.B(\macro_inst|ahb_add_reg [18]),
	.C(\rv32.mem_ahb_haddr[17] ),
	.D(\macro_inst|ahb_add_reg [19]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [17]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X57_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y3_SIG ),
	.SyncReset(SyncReset_X57_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|motor_flags[0]~4_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [17]));
defparam \macro_inst|ahb_add_reg[17] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[17] .coord_y = 11;
defparam \macro_inst|ahb_add_reg[17] .coord_z = 1;
defparam \macro_inst|ahb_add_reg[17] .mask = 16'h0001;
defparam \macro_inst|ahb_add_reg[17] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[17] .FeedbackMux = 1'b1;
defparam \macro_inst|ahb_add_reg[17] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[17] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[17] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[18] (
	.A(\rv32.mem_ahb_haddr[31] ),
	.B(\rv32.mem_ahb_haddr[27] ),
	.C(\rv32.mem_ahb_haddr[18] ),
	.D(\rv32.mem_ahb_haddr[17] ),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [18]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X57_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y3_SIG ),
	.SyncReset(SyncReset_X57_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y3_VCC),
	.LutOut(\macro_inst|Equal1~5_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [18]));
defparam \macro_inst|ahb_add_reg[18] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[18] .coord_y = 11;
defparam \macro_inst|ahb_add_reg[18] .coord_z = 13;
defparam \macro_inst|ahb_add_reg[18] .mask = 16'h0001;
defparam \macro_inst|ahb_add_reg[18] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[18] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[18] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[18] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[18] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[19] (
	.A(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [19]),
	.B(vcc),
	.C(\rv32.mem_ahb_haddr[19] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [19]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X57_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y3_SIG ),
	.SyncReset(SyncReset_X57_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y3_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[19]~19_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [19]));
defparam \macro_inst|ahb_add_reg[19] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[19] .coord_y = 11;
defparam \macro_inst|ahb_add_reg[19] .coord_z = 3;
defparam \macro_inst|ahb_add_reg[19] .mask = 16'hAA00;
defparam \macro_inst|ahb_add_reg[19] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[19] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[19] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[19] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[19] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[1] (
	.A(\macro_inst|ahb_add_reg [3]),
	.B(vcc),
	.C(\rv32.mem_ahb_haddr[1] ),
	.D(\macro_inst|ahb_add_reg [2]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X60_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y3_SIG ),
	.SyncReset(SyncReset_X60_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~18_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [1]));
defparam \macro_inst|ahb_add_reg[1] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[1] .coord_y = 7;
defparam \macro_inst|ahb_add_reg[1] .coord_z = 5;
defparam \macro_inst|ahb_add_reg[1] .mask = 16'hAA00;
defparam \macro_inst|ahb_add_reg[1] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[1] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[1] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[1] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[1] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[20] (
	.A(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [20]),
	.B(vcc),
	.C(\rv32.mem_ahb_haddr[20] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [20]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X57_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y3_SIG ),
	.SyncReset(SyncReset_X57_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y3_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[20]~20_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [20]));
defparam \macro_inst|ahb_add_reg[20] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[20] .coord_y = 11;
defparam \macro_inst|ahb_add_reg[20] .coord_z = 8;
defparam \macro_inst|ahb_add_reg[20] .mask = 16'hAA00;
defparam \macro_inst|ahb_add_reg[20] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[20] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[20] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[20] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[20] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[21] (
	.A(\macro_inst|ahb_add_reg [22]),
	.B(\macro_inst|ahb_add_reg [24]),
	.C(\rv32.mem_ahb_haddr[21] ),
	.D(\macro_inst|ahb_add_reg [23]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [21]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(SyncReset_X54_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|motor_flags[0]~2_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [21]));
defparam \macro_inst|ahb_add_reg[21] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[21] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[21] .coord_z = 6;
defparam \macro_inst|ahb_add_reg[21] .mask = 16'h0001;
defparam \macro_inst|ahb_add_reg[21] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[21] .FeedbackMux = 1'b1;
defparam \macro_inst|ahb_add_reg[21] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[21] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[21] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[22] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [22]),
	.C(\rv32.mem_ahb_haddr[22] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [22]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(SyncReset_X54_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y3_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[22]~22_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [22]));
defparam \macro_inst|ahb_add_reg[22] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[22] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[22] .coord_z = 0;
defparam \macro_inst|ahb_add_reg[22] .mask = 16'hCC00;
defparam \macro_inst|ahb_add_reg[22] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[22] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[22] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[22] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[22] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[23] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [23]),
	.C(\rv32.mem_ahb_haddr[23] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [23]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(SyncReset_X54_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y3_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[23]~23_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [23]));
defparam \macro_inst|ahb_add_reg[23] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[23] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[23] .coord_z = 11;
defparam \macro_inst|ahb_add_reg[23] .mask = 16'hCC00;
defparam \macro_inst|ahb_add_reg[23] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[23] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[23] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[23] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[23] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[24] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [24]),
	.C(\rv32.mem_ahb_haddr[24] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [24]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(SyncReset_X54_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y3_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[24]~24_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [24]));
defparam \macro_inst|ahb_add_reg[24] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[24] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[24] .coord_z = 1;
defparam \macro_inst|ahb_add_reg[24] .mask = 16'hCC00;
defparam \macro_inst|ahb_add_reg[24] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[24] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[24] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[24] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[24] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[25] (
	.A(\macro_inst|ahb_add_reg [28]),
	.B(\macro_inst|ahb_add_reg [27]),
	.C(\rv32.mem_ahb_haddr[25] ),
	.D(\macro_inst|ahb_add_reg [26]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [25]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(SyncReset_X54_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|motor_flags[0]~1_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [25]));
defparam \macro_inst|ahb_add_reg[25] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[25] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[25] .coord_z = 12;
defparam \macro_inst|ahb_add_reg[25] .mask = 16'h0001;
defparam \macro_inst|ahb_add_reg[25] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[25] .FeedbackMux = 1'b1;
defparam \macro_inst|ahb_add_reg[25] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[25] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[25] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[26] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [26]),
	.C(\rv32.mem_ahb_haddr[26] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [26]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(SyncReset_X54_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y3_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[26]~26_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [26]));
defparam \macro_inst|ahb_add_reg[26] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[26] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[26] .coord_z = 3;
defparam \macro_inst|ahb_add_reg[26] .mask = 16'hCC00;
defparam \macro_inst|ahb_add_reg[26] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[26] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[26] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[26] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[26] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[27] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [27]),
	.C(\rv32.mem_ahb_haddr[27] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [27]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(SyncReset_X54_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y3_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[27]~27_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [27]));
defparam \macro_inst|ahb_add_reg[27] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[27] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[27] .coord_z = 15;
defparam \macro_inst|ahb_add_reg[27] .mask = 16'hCC00;
defparam \macro_inst|ahb_add_reg[27] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[27] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[27] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[27] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[27] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[28] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [28]),
	.C(\rv32.mem_ahb_haddr[28] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [28]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(SyncReset_X54_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y3_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[28]~28_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [28]));
defparam \macro_inst|ahb_add_reg[28] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[28] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[28] .coord_z = 4;
defparam \macro_inst|ahb_add_reg[28] .mask = 16'hCC00;
defparam \macro_inst|ahb_add_reg[28] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[28] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[28] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[28] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[28] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[29] (
	.A(\macro_inst|ahb_ready_reg~q ),
	.B(\macro_inst|ahb_add_reg [31]),
	.C(\rv32.mem_ahb_haddr[29] ),
	.D(\macro_inst|ahb_add_reg [30]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [29]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X57_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y3_SIG ),
	.SyncReset(SyncReset_X57_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|motor_flags[0]~0_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [29]));
defparam \macro_inst|ahb_add_reg[29] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[29] .coord_y = 11;
defparam \macro_inst|ahb_add_reg[29] .coord_z = 11;
defparam \macro_inst|ahb_add_reg[29] .mask = 16'h2000;
defparam \macro_inst|ahb_add_reg[29] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[29] .FeedbackMux = 1'b1;
defparam \macro_inst|ahb_add_reg[29] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[29] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[29] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[2] (
	.A(\macro_inst|ahb_add_reg [4]),
	.B(\macro_inst|ahb_add_reg [5]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|ahb_add_reg [1]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X60_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y3_SIG ),
	.SyncReset(SyncReset_X60_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~13_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [2]));
defparam \macro_inst|ahb_add_reg[2] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[2] .coord_y = 7;
defparam \macro_inst|ahb_add_reg[2] .coord_z = 11;
defparam \macro_inst|ahb_add_reg[2] .mask = 16'h1100;
defparam \macro_inst|ahb_add_reg[2] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[2] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[2] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[2] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[2] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[30] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [30]),
	.C(\rv32.mem_ahb_haddr[30] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [30]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X57_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y3_SIG ),
	.SyncReset(SyncReset_X57_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y3_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[30]~30_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [30]));
defparam \macro_inst|ahb_add_reg[30] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[30] .coord_y = 11;
defparam \macro_inst|ahb_add_reg[30] .coord_z = 15;
defparam \macro_inst|ahb_add_reg[30] .mask = 16'hCC00;
defparam \macro_inst|ahb_add_reg[30] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[30] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[30] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[30] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[30] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[31] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [31]),
	.C(\rv32.mem_ahb_haddr[31] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [31]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X57_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y3_SIG ),
	.SyncReset(SyncReset_X57_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y3_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[31]~31_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [31]));
defparam \macro_inst|ahb_add_reg[31] .coord_x = 14;
defparam \macro_inst|ahb_add_reg[31] .coord_y = 11;
defparam \macro_inst|ahb_add_reg[31] .coord_z = 5;
defparam \macro_inst|ahb_add_reg[31] .mask = 16'hCC00;
defparam \macro_inst|ahb_add_reg[31] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[31] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[31] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[31] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[31] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[3] (
	.A(vcc),
	.B(vcc),
	.C(\rv32.mem_ahb_haddr[3] ),
	.D(\macro_inst|ahb_add_reg [2]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [3]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X60_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y3_SIG ),
	.SyncReset(SyncReset_X60_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~4_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [3]));
defparam \macro_inst|ahb_add_reg[3] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[3] .coord_y = 7;
defparam \macro_inst|ahb_add_reg[3] .coord_z = 6;
defparam \macro_inst|ahb_add_reg[3] .mask = 16'h000F;
defparam \macro_inst|ahb_add_reg[3] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[3] .FeedbackMux = 1'b1;
defparam \macro_inst|ahb_add_reg[3] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[3] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[3] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[4] (
	.A(vcc),
	.B(\macro_inst|ahb_add_reg [6]),
	.C(\rv32.mem_ahb_haddr[4] ),
	.D(\macro_inst|ahb_add_reg [5]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [4]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X60_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y3_SIG ),
	.SyncReset(SyncReset_X60_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~35_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [4]));
defparam \macro_inst|ahb_add_reg[4] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[4] .coord_y = 7;
defparam \macro_inst|ahb_add_reg[4] .coord_z = 14;
defparam \macro_inst|ahb_add_reg[4] .mask = 16'h00C0;
defparam \macro_inst|ahb_add_reg[4] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[4] .FeedbackMux = 1'b1;
defparam \macro_inst|ahb_add_reg[4] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[4] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[4] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[5] (
	.A(\macro_inst|ahb_add_reg [4]),
	.B(vcc),
	.C(\rv32.mem_ahb_haddr[5] ),
	.D(\macro_inst|ahb_add_reg [6]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [5]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X58_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y3_SIG ),
	.SyncReset(SyncReset_X58_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~75_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [5]));
defparam \macro_inst|ahb_add_reg[5] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[5] .coord_y = 11;
defparam \macro_inst|ahb_add_reg[5] .coord_z = 1;
defparam \macro_inst|ahb_add_reg[5] .mask = 16'h000A;
defparam \macro_inst|ahb_add_reg[5] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[5] .FeedbackMux = 1'b1;
defparam \macro_inst|ahb_add_reg[5] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[5] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[5] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[6] (
	.A(\macro_inst|controller|sm_pwm|Decoder0~13_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~12_combout ),
	.C(\rv32.mem_ahb_haddr[6] ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [6]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X59_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y3_SIG ),
	.SyncReset(SyncReset_X59_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~14_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [6]));
defparam \macro_inst|ahb_add_reg[6] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[6] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[6] .coord_z = 14;
defparam \macro_inst|ahb_add_reg[6] .mask = 16'h0800;
defparam \macro_inst|ahb_add_reg[6] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[6] .FeedbackMux = 1'b1;
defparam \macro_inst|ahb_add_reg[6] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[6] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[6] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[7] (
	.A(\macro_inst|ahb_add_reg [6]),
	.B(\macro_inst|ahb_add_reg [5]),
	.C(\rv32.mem_ahb_haddr[7] ),
	.D(\macro_inst|ahb_add_reg [1]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [7]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X59_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y3_SIG ),
	.SyncReset(SyncReset_X59_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~53_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [7]));
defparam \macro_inst|ahb_add_reg[7] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[7] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[7] .coord_z = 15;
defparam \macro_inst|ahb_add_reg[7] .mask = 16'h0044;
defparam \macro_inst|ahb_add_reg[7] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[7] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[7] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[7] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[7] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[8] (
	.A(\macro_inst|ahb_add_reg [10]),
	.B(\macro_inst|ahb_add_reg [9]),
	.C(\rv32.mem_ahb_haddr[8] ),
	.D(\macro_inst|ahb_add_reg [11]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [8]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X59_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y3_SIG ),
	.SyncReset(SyncReset_X59_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~7_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [8]));
defparam \macro_inst|ahb_add_reg[8] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[8] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[8] .coord_z = 1;
defparam \macro_inst|ahb_add_reg[8] .mask = 16'h0001;
defparam \macro_inst|ahb_add_reg[8] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[8] .FeedbackMux = 1'b1;
defparam \macro_inst|ahb_add_reg[8] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[8] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[8] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_add_reg[9] (
	.A(\macro_inst|ahb_add_reg [6]),
	.B(\macro_inst|ahb_add_reg [5]),
	.C(\rv32.mem_ahb_haddr[9] ),
	.D(\macro_inst|ahb_add_reg [1]),
	.Cin(),
	.Qin(\macro_inst|ahb_add_reg [9]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X59_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y3_SIG ),
	.SyncReset(SyncReset_X59_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~71_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_add_reg [9]));
defparam \macro_inst|ahb_add_reg[9] .coord_x = 15;
defparam \macro_inst|ahb_add_reg[9] .coord_y = 12;
defparam \macro_inst|ahb_add_reg[9] .coord_z = 0;
defparam \macro_inst|ahb_add_reg[9] .mask = 16'h0011;
defparam \macro_inst|ahb_add_reg[9] .modeMux = 1'b0;
defparam \macro_inst|ahb_add_reg[9] .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_add_reg[9] .ShiftMux = 1'b0;
defparam \macro_inst|ahb_add_reg[9] .BypassEn = 1'b1;
defparam \macro_inst|ahb_add_reg[9] .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_ready_reg (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [29]),
	.C(\macro_inst|Equal2~0_combout ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_ready_reg~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y3_SIG ),
	.SyncReset(SyncReset_X57_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y3_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[29]~29_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_ready_reg~q ));
defparam \macro_inst|ahb_ready_reg .coord_x = 14;
defparam \macro_inst|ahb_ready_reg .coord_y = 11;
defparam \macro_inst|ahb_ready_reg .coord_z = 4;
defparam \macro_inst|ahb_ready_reg .mask = 16'hCC00;
defparam \macro_inst|ahb_ready_reg .modeMux = 1'b0;
defparam \macro_inst|ahb_ready_reg .FeedbackMux = 1'b0;
defparam \macro_inst|ahb_ready_reg .ShiftMux = 1'b0;
defparam \macro_inst|ahb_ready_reg .BypassEn = 1'b1;
defparam \macro_inst|ahb_ready_reg .CarryEnb = 1'b1;

alta_slice \macro_inst|ahb_wr_reg (
	.A(\macro_inst|ahb_add_reg [16]),
	.B(vcc),
	.C(\rv32.mem_ahb_hwrite ),
	.D(\macro_inst|controller|sm_pwm|motor_flags[0]~4_combout ),
	.Cin(),
	.Qin(\macro_inst|ahb_wr_reg~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|Equal2~0_combout_X58_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y3_SIG ),
	.SyncReset(SyncReset_X58_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|motor_flags[0]~5_combout ),
	.Cout(),
	.Q(\macro_inst|ahb_wr_reg~q ));
defparam \macro_inst|ahb_wr_reg .coord_x = 15;
defparam \macro_inst|ahb_wr_reg .coord_y = 11;
defparam \macro_inst|ahb_wr_reg .coord_z = 11;
defparam \macro_inst|ahb_wr_reg .mask = 16'h5000;
defparam \macro_inst|ahb_wr_reg .modeMux = 1'b0;
defparam \macro_inst|ahb_wr_reg .FeedbackMux = 1'b1;
defparam \macro_inst|ahb_wr_reg .ShiftMux = 1'b0;
defparam \macro_inst|ahb_wr_reg .BypassEn = 1'b1;
defparam \macro_inst|ahb_wr_reg .CarryEnb = 1'b1;

alta_slice \macro_inst|clk10hz_cnt[0] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|clk10hz_cnt [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~0_combout ),
	.Cout(\macro_inst|Add0~1 ),
	.Q(\macro_inst|clk10hz_cnt [0]));
defparam \macro_inst|clk10hz_cnt[0] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[0] .coord_y = 2;
defparam \macro_inst|clk10hz_cnt[0] .coord_z = 5;
defparam \macro_inst|clk10hz_cnt[0] .mask = 16'h33CC;
defparam \macro_inst|clk10hz_cnt[0] .modeMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[0] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[0] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[0] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[0] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[10] (
	.A(\macro_inst|Equal3~5_combout ),
	.B(\macro_inst|Add0~20_combout ),
	.C(\macro_inst|Equal3~4_combout ),
	.D(\macro_inst|Equal3~6_combout ),
	.Cin(),
	.Qin(\macro_inst|clk10hz_cnt [10]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|clk10hz_cnt~1_combout ),
	.Cout(),
	.Q(\macro_inst|clk10hz_cnt [10]));
defparam \macro_inst|clk10hz_cnt[10] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[10] .coord_y = 2;
defparam \macro_inst|clk10hz_cnt[10] .coord_z = 4;
defparam \macro_inst|clk10hz_cnt[10] .mask = 16'h4CCC;
defparam \macro_inst|clk10hz_cnt[10] .modeMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[10] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[10] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[10] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[10] .CarryEnb = 1'b1;

alta_slice \macro_inst|clk10hz_cnt[11] (
	.A(\macro_inst|Add0~22_combout ),
	.B(\macro_inst|Equal3~5_combout ),
	.C(\macro_inst|Equal3~6_combout ),
	.D(\macro_inst|Equal3~4_combout ),
	.Cin(),
	.Qin(\macro_inst|clk10hz_cnt [11]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X47_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X47_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|clk10hz_cnt~0_combout ),
	.Cout(),
	.Q(\macro_inst|clk10hz_cnt [11]));
defparam \macro_inst|clk10hz_cnt[11] .coord_x = 4;
defparam \macro_inst|clk10hz_cnt[11] .coord_y = 2;
defparam \macro_inst|clk10hz_cnt[11] .coord_z = 7;
defparam \macro_inst|clk10hz_cnt[11] .mask = 16'h2AAA;
defparam \macro_inst|clk10hz_cnt[11] .modeMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[11] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[11] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[11] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[11] .CarryEnb = 1'b1;

alta_slice \macro_inst|clk10hz_cnt[12] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [12]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~23 ),
	.Qin(\macro_inst|clk10hz_cnt [12]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~24_combout ),
	.Cout(\macro_inst|Add0~25 ),
	.Q(\macro_inst|clk10hz_cnt [12]));
defparam \macro_inst|clk10hz_cnt[12] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[12] .coord_y = 1;
defparam \macro_inst|clk10hz_cnt[12] .coord_z = 1;
defparam \macro_inst|clk10hz_cnt[12] .mask = 16'hC30C;
defparam \macro_inst|clk10hz_cnt[12] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[12] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[12] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[12] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[12] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[13] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [13]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~25 ),
	.Qin(\macro_inst|clk10hz_cnt [13]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~26_combout ),
	.Cout(\macro_inst|Add0~27 ),
	.Q(\macro_inst|clk10hz_cnt [13]));
defparam \macro_inst|clk10hz_cnt[13] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[13] .coord_y = 1;
defparam \macro_inst|clk10hz_cnt[13] .coord_z = 2;
defparam \macro_inst|clk10hz_cnt[13] .mask = 16'h3C3F;
defparam \macro_inst|clk10hz_cnt[13] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[13] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[13] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[13] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[13] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[14] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [14]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~27 ),
	.Qin(\macro_inst|clk10hz_cnt [14]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~28_combout ),
	.Cout(\macro_inst|Add0~29 ),
	.Q(\macro_inst|clk10hz_cnt [14]));
defparam \macro_inst|clk10hz_cnt[14] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[14] .coord_y = 1;
defparam \macro_inst|clk10hz_cnt[14] .coord_z = 3;
defparam \macro_inst|clk10hz_cnt[14] .mask = 16'hC30C;
defparam \macro_inst|clk10hz_cnt[14] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[14] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[14] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[14] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[14] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[15] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [15]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~29 ),
	.Qin(\macro_inst|clk10hz_cnt [15]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~30_combout ),
	.Cout(\macro_inst|Add0~31 ),
	.Q(\macro_inst|clk10hz_cnt [15]));
defparam \macro_inst|clk10hz_cnt[15] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[15] .coord_y = 1;
defparam \macro_inst|clk10hz_cnt[15] .coord_z = 4;
defparam \macro_inst|clk10hz_cnt[15] .mask = 16'h3C3F;
defparam \macro_inst|clk10hz_cnt[15] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[15] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[15] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[15] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[15] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[16] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [16]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~31 ),
	.Qin(\macro_inst|clk10hz_cnt [16]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~32_combout ),
	.Cout(\macro_inst|Add0~33 ),
	.Q(\macro_inst|clk10hz_cnt [16]));
defparam \macro_inst|clk10hz_cnt[16] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[16] .coord_y = 1;
defparam \macro_inst|clk10hz_cnt[16] .coord_z = 5;
defparam \macro_inst|clk10hz_cnt[16] .mask = 16'hC30C;
defparam \macro_inst|clk10hz_cnt[16] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[16] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[16] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[16] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[16] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[17] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [17]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~33 ),
	.Qin(\macro_inst|clk10hz_cnt [17]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~34_combout ),
	.Cout(\macro_inst|Add0~35 ),
	.Q(\macro_inst|clk10hz_cnt [17]));
defparam \macro_inst|clk10hz_cnt[17] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[17] .coord_y = 1;
defparam \macro_inst|clk10hz_cnt[17] .coord_z = 6;
defparam \macro_inst|clk10hz_cnt[17] .mask = 16'h3C3F;
defparam \macro_inst|clk10hz_cnt[17] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[17] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[17] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[17] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[17] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[18] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [18]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~35 ),
	.Qin(\macro_inst|clk10hz_cnt [18]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~36_combout ),
	.Cout(\macro_inst|Add0~37 ),
	.Q(\macro_inst|clk10hz_cnt [18]));
defparam \macro_inst|clk10hz_cnt[18] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[18] .coord_y = 1;
defparam \macro_inst|clk10hz_cnt[18] .coord_z = 7;
defparam \macro_inst|clk10hz_cnt[18] .mask = 16'hC30C;
defparam \macro_inst|clk10hz_cnt[18] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[18] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[18] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[18] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[18] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[19] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [19]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~37 ),
	.Qin(\macro_inst|clk10hz_cnt [19]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~38_combout ),
	.Cout(\macro_inst|Add0~39 ),
	.Q(\macro_inst|clk10hz_cnt [19]));
defparam \macro_inst|clk10hz_cnt[19] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[19] .coord_y = 1;
defparam \macro_inst|clk10hz_cnt[19] .coord_z = 8;
defparam \macro_inst|clk10hz_cnt[19] .mask = 16'h3C3F;
defparam \macro_inst|clk10hz_cnt[19] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[19] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[19] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[19] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[19] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[1] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~1 ),
	.Qin(\macro_inst|clk10hz_cnt [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~2_combout ),
	.Cout(\macro_inst|Add0~3 ),
	.Q(\macro_inst|clk10hz_cnt [1]));
defparam \macro_inst|clk10hz_cnt[1] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[1] .coord_y = 2;
defparam \macro_inst|clk10hz_cnt[1] .coord_z = 6;
defparam \macro_inst|clk10hz_cnt[1] .mask = 16'h3C3F;
defparam \macro_inst|clk10hz_cnt[1] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[1] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[1] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[1] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[1] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[20] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [20]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~39 ),
	.Qin(\macro_inst|clk10hz_cnt [20]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~40_combout ),
	.Cout(\macro_inst|Add0~41 ),
	.Q(\macro_inst|clk10hz_cnt [20]));
defparam \macro_inst|clk10hz_cnt[20] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[20] .coord_y = 1;
defparam \macro_inst|clk10hz_cnt[20] .coord_z = 9;
defparam \macro_inst|clk10hz_cnt[20] .mask = 16'hC30C;
defparam \macro_inst|clk10hz_cnt[20] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[20] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[20] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[20] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[20] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[21] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [21]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~41 ),
	.Qin(\macro_inst|clk10hz_cnt [21]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~42_combout ),
	.Cout(\macro_inst|Add0~43 ),
	.Q(\macro_inst|clk10hz_cnt [21]));
defparam \macro_inst|clk10hz_cnt[21] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[21] .coord_y = 1;
defparam \macro_inst|clk10hz_cnt[21] .coord_z = 10;
defparam \macro_inst|clk10hz_cnt[21] .mask = 16'h3C3F;
defparam \macro_inst|clk10hz_cnt[21] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[21] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[21] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[21] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[21] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[22] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [22]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~43 ),
	.Qin(\macro_inst|clk10hz_cnt [22]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~44_combout ),
	.Cout(),
	.Q(\macro_inst|clk10hz_cnt [22]));
defparam \macro_inst|clk10hz_cnt[22] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[22] .coord_y = 1;
defparam \macro_inst|clk10hz_cnt[22] .coord_z = 11;
defparam \macro_inst|clk10hz_cnt[22] .mask = 16'hC3C3;
defparam \macro_inst|clk10hz_cnt[22] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[22] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[22] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[22] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[22] .CarryEnb = 1'b1;

alta_slice \macro_inst|clk10hz_cnt[2] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~3 ),
	.Qin(\macro_inst|clk10hz_cnt [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~4_combout ),
	.Cout(\macro_inst|Add0~5 ),
	.Q(\macro_inst|clk10hz_cnt [2]));
defparam \macro_inst|clk10hz_cnt[2] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[2] .coord_y = 2;
defparam \macro_inst|clk10hz_cnt[2] .coord_z = 7;
defparam \macro_inst|clk10hz_cnt[2] .mask = 16'hC30C;
defparam \macro_inst|clk10hz_cnt[2] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[2] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[2] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[2] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[2] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[3] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~5 ),
	.Qin(\macro_inst|clk10hz_cnt [3]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~6_combout ),
	.Cout(\macro_inst|Add0~7 ),
	.Q(\macro_inst|clk10hz_cnt [3]));
defparam \macro_inst|clk10hz_cnt[3] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[3] .coord_y = 2;
defparam \macro_inst|clk10hz_cnt[3] .coord_z = 8;
defparam \macro_inst|clk10hz_cnt[3] .mask = 16'h3C3F;
defparam \macro_inst|clk10hz_cnt[3] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[3] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[3] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[3] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[3] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[4] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~7 ),
	.Qin(\macro_inst|clk10hz_cnt [4]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~8_combout ),
	.Cout(\macro_inst|Add0~9 ),
	.Q(\macro_inst|clk10hz_cnt [4]));
defparam \macro_inst|clk10hz_cnt[4] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[4] .coord_y = 2;
defparam \macro_inst|clk10hz_cnt[4] .coord_z = 9;
defparam \macro_inst|clk10hz_cnt[4] .mask = 16'hC30C;
defparam \macro_inst|clk10hz_cnt[4] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[4] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[4] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[4] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[4] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[5] (
	.A(\macro_inst|Add0~10_combout ),
	.B(\macro_inst|Equal3~6_combout ),
	.C(\macro_inst|Equal3~5_combout ),
	.D(\macro_inst|Equal3~4_combout ),
	.Cin(),
	.Qin(\macro_inst|clk10hz_cnt [5]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|clk10hz_cnt~5_combout ),
	.Cout(),
	.Q(\macro_inst|clk10hz_cnt [5]));
defparam \macro_inst|clk10hz_cnt[5] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[5] .coord_y = 2;
defparam \macro_inst|clk10hz_cnt[5] .coord_z = 1;
defparam \macro_inst|clk10hz_cnt[5] .mask = 16'h2AAA;
defparam \macro_inst|clk10hz_cnt[5] .modeMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[5] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[5] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[5] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[5] .CarryEnb = 1'b1;

alta_slice \macro_inst|clk10hz_cnt[6] (
	.A(vcc),
	.B(\macro_inst|clk10hz_cnt [6]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|Add0~11 ),
	.Qin(\macro_inst|clk10hz_cnt [6]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|Add0~12_combout ),
	.Cout(\macro_inst|Add0~13 ),
	.Q(\macro_inst|clk10hz_cnt [6]));
defparam \macro_inst|clk10hz_cnt[6] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[6] .coord_y = 2;
defparam \macro_inst|clk10hz_cnt[6] .coord_z = 11;
defparam \macro_inst|clk10hz_cnt[6] .mask = 16'hC30C;
defparam \macro_inst|clk10hz_cnt[6] .modeMux = 1'b1;
defparam \macro_inst|clk10hz_cnt[6] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[6] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[6] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[6] .CarryEnb = 1'b0;

alta_slice \macro_inst|clk10hz_cnt[7] (
	.A(\macro_inst|Add0~14_combout ),
	.B(\macro_inst|Equal3~5_combout ),
	.C(\macro_inst|Equal3~6_combout ),
	.D(\macro_inst|Equal3~4_combout ),
	.Cin(),
	.Qin(\macro_inst|clk10hz_cnt [7]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X47_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X47_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|clk10hz_cnt~4_combout ),
	.Cout(),
	.Q(\macro_inst|clk10hz_cnt [7]));
defparam \macro_inst|clk10hz_cnt[7] .coord_x = 4;
defparam \macro_inst|clk10hz_cnt[7] .coord_y = 2;
defparam \macro_inst|clk10hz_cnt[7] .coord_z = 5;
defparam \macro_inst|clk10hz_cnt[7] .mask = 16'h2AAA;
defparam \macro_inst|clk10hz_cnt[7] .modeMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[7] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[7] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[7] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[7] .CarryEnb = 1'b1;

alta_slice \macro_inst|clk10hz_cnt[8] (
	.A(\macro_inst|Equal3~5_combout ),
	.B(\macro_inst|Add0~16_combout ),
	.C(\macro_inst|Equal3~4_combout ),
	.D(\macro_inst|Equal3~6_combout ),
	.Cin(),
	.Qin(\macro_inst|clk10hz_cnt [8]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|clk10hz_cnt~3_combout ),
	.Cout(),
	.Q(\macro_inst|clk10hz_cnt [8]));
defparam \macro_inst|clk10hz_cnt[8] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[8] .coord_y = 2;
defparam \macro_inst|clk10hz_cnt[8] .coord_z = 0;
defparam \macro_inst|clk10hz_cnt[8] .mask = 16'h4CCC;
defparam \macro_inst|clk10hz_cnt[8] .modeMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[8] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[8] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[8] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[8] .CarryEnb = 1'b1;

alta_slice \macro_inst|clk10hz_cnt[9] (
	.A(\macro_inst|Add0~18_combout ),
	.B(\macro_inst|Equal3~6_combout ),
	.C(\macro_inst|Equal3~5_combout ),
	.D(\macro_inst|Equal3~4_combout ),
	.Cin(),
	.Qin(\macro_inst|clk10hz_cnt [9]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X48_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X48_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|clk10hz_cnt~2_combout ),
	.Cout(),
	.Q(\macro_inst|clk10hz_cnt [9]));
defparam \macro_inst|clk10hz_cnt[9] .coord_x = 3;
defparam \macro_inst|clk10hz_cnt[9] .coord_y = 2;
defparam \macro_inst|clk10hz_cnt[9] .coord_z = 3;
defparam \macro_inst|clk10hz_cnt[9] .mask = 16'h2AAA;
defparam \macro_inst|clk10hz_cnt[9] .modeMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[9] .FeedbackMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[9] .ShiftMux = 1'b0;
defparam \macro_inst|clk10hz_cnt[9] .BypassEn = 1'b0;
defparam \macro_inst|clk10hz_cnt[9] .CarryEnb = 1'b1;

alta_slice \macro_inst|clock10Hz (
	.A(\macro_inst|Equal3~6_combout ),
	.B(\macro_inst|Equal3~5_combout ),
	.C(vcc),
	.D(\macro_inst|Equal3~4_combout ),
	.Cin(),
	.Qin(\macro_inst|clock10Hz~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X47_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X47_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|clock10Hz~0_combout ),
	.Cout(),
	.Q(\macro_inst|clock10Hz~q ));
defparam \macro_inst|clock10Hz .coord_x = 4;
defparam \macro_inst|clock10Hz .coord_y = 2;
defparam \macro_inst|clock10Hz .coord_z = 8;
defparam \macro_inst|clock10Hz .mask = 16'h78F0;
defparam \macro_inst|clock10Hz .modeMux = 1'b0;
defparam \macro_inst|clock10Hz .FeedbackMux = 1'b1;
defparam \macro_inst|clock10Hz .ShiftMux = 1'b0;
defparam \macro_inst|clock10Hz .BypassEn = 1'b0;
defparam \macro_inst|clock10Hz .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|Add0~0 (
	.A(\macro_inst|controller|serialTrigCounter [0]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|Add0~0_combout ),
	.Cout(\macro_inst|controller|Add0~1 ),
	.Q());
defparam \macro_inst|controller|Add0~0 .coord_x = 6;
defparam \macro_inst|controller|Add0~0 .coord_y = 1;
defparam \macro_inst|controller|Add0~0 .coord_z = 5;
defparam \macro_inst|controller|Add0~0 .mask = 16'h55AA;
defparam \macro_inst|controller|Add0~0 .modeMux = 1'b0;
defparam \macro_inst|controller|Add0~0 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|Add0~0 .ShiftMux = 1'b0;
defparam \macro_inst|controller|Add0~0 .BypassEn = 1'b0;
defparam \macro_inst|controller|Add0~0 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|Add0~10 (
	.A(vcc),
	.B(\macro_inst|controller|serialTrigCounter [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|Add0~9 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|Add0~10_combout ),
	.Cout(\macro_inst|controller|Add0~11 ),
	.Q());
defparam \macro_inst|controller|Add0~10 .coord_x = 6;
defparam \macro_inst|controller|Add0~10 .coord_y = 1;
defparam \macro_inst|controller|Add0~10 .coord_z = 10;
defparam \macro_inst|controller|Add0~10 .mask = 16'h3C3F;
defparam \macro_inst|controller|Add0~10 .modeMux = 1'b1;
defparam \macro_inst|controller|Add0~10 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|Add0~10 .ShiftMux = 1'b0;
defparam \macro_inst|controller|Add0~10 .BypassEn = 1'b0;
defparam \macro_inst|controller|Add0~10 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|Add0~4 (
	.A(vcc),
	.B(\macro_inst|controller|serialTrigCounter [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|Add0~3 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|Add0~4_combout ),
	.Cout(\macro_inst|controller|Add0~5 ),
	.Q());
defparam \macro_inst|controller|Add0~4 .coord_x = 6;
defparam \macro_inst|controller|Add0~4 .coord_y = 1;
defparam \macro_inst|controller|Add0~4 .coord_z = 7;
defparam \macro_inst|controller|Add0~4 .mask = 16'hC30C;
defparam \macro_inst|controller|Add0~4 .modeMux = 1'b1;
defparam \macro_inst|controller|Add0~4 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|Add0~4 .ShiftMux = 1'b0;
defparam \macro_inst|controller|Add0~4 .BypassEn = 1'b0;
defparam \macro_inst|controller|Add0~4 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|Equal1~0 (
	.A(\macro_inst|controller|serialTrigCounter [6]),
	.B(\macro_inst|controller|serialTrigCounter [5]),
	.C(\macro_inst|controller|serialTrigCounter [7]),
	.D(\macro_inst|controller|serialTrigCounter [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|Equal1~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|Equal1~0 .coord_x = 6;
defparam \macro_inst|controller|Equal1~0 .coord_y = 1;
defparam \macro_inst|controller|Equal1~0 .coord_z = 0;
defparam \macro_inst|controller|Equal1~0 .mask = 16'h0004;
defparam \macro_inst|controller|Equal1~0 .modeMux = 1'b0;
defparam \macro_inst|controller|Equal1~0 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|Equal1~0 .ShiftMux = 1'b0;
defparam \macro_inst|controller|Equal1~0 .BypassEn = 1'b0;
defparam \macro_inst|controller|Equal1~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|Equal1~1 (
	.A(\macro_inst|controller|serialTrigCounter [1]),
	.B(\macro_inst|controller|serialTrigCounter [3]),
	.C(\macro_inst|controller|serialTrigCounter [0]),
	.D(\macro_inst|controller|serialTrigCounter [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|Equal1~1_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|Equal1~1 .coord_x = 6;
defparam \macro_inst|controller|Equal1~1 .coord_y = 1;
defparam \macro_inst|controller|Equal1~1 .coord_z = 14;
defparam \macro_inst|controller|Equal1~1 .mask = 16'h0100;
defparam \macro_inst|controller|Equal1~1 .modeMux = 1'b0;
defparam \macro_inst|controller|Equal1~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|Equal1~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|Equal1~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|Equal1~1 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|Equal1~2 (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|Equal1~0_combout ),
	.D(\macro_inst|controller|Equal1~1_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|Equal1~2_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|Equal1~2 .coord_x = 7;
defparam \macro_inst|controller|Equal1~2 .coord_y = 1;
defparam \macro_inst|controller|Equal1~2 .coord_z = 0;
defparam \macro_inst|controller|Equal1~2 .mask = 16'hF000;
defparam \macro_inst|controller|Equal1~2 .modeMux = 1'b0;
defparam \macro_inst|controller|Equal1~2 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|Equal1~2 .ShiftMux = 1'b0;
defparam \macro_inst|controller|Equal1~2 .BypassEn = 1'b0;
defparam \macro_inst|controller|Equal1~2 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|pwmUpdateTrigger (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|Equal1~2_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|pwmUpdateTrigger~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X51_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|pwmUpdateTrigger~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|pwmUpdateTrigger~q ));
defparam \macro_inst|controller|pwmUpdateTrigger .coord_x = 8;
defparam \macro_inst|controller|pwmUpdateTrigger .coord_y = 1;
defparam \macro_inst|controller|pwmUpdateTrigger .coord_z = 1;
defparam \macro_inst|controller|pwmUpdateTrigger .mask = 16'hFF00;
defparam \macro_inst|controller|pwmUpdateTrigger .modeMux = 1'b0;
defparam \macro_inst|controller|pwmUpdateTrigger .FeedbackMux = 1'b0;
defparam \macro_inst|controller|pwmUpdateTrigger .ShiftMux = 1'b0;
defparam \macro_inst|controller|pwmUpdateTrigger .BypassEn = 1'b0;
defparam \macro_inst|controller|pwmUpdateTrigger .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serialOutputTrigger[0] (
	.A(\macro_inst|controller|serialOutputTrigger [1]),
	.B(\macro_inst|controller|pwmUpdateTrigger~q ),
	.C(vcc),
	.D(\macro_inst|controller|Equal1~2_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serialOutputTrigger [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X51_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serialOutputTrigger[0]~1_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serialOutputTrigger [0]));
defparam \macro_inst|controller|serialOutputTrigger[0] .coord_x = 8;
defparam \macro_inst|controller|serialOutputTrigger[0] .coord_y = 1;
defparam \macro_inst|controller|serialOutputTrigger[0] .coord_z = 13;
defparam \macro_inst|controller|serialOutputTrigger[0] .mask = 16'hF002;
defparam \macro_inst|controller|serialOutputTrigger[0] .modeMux = 1'b0;
defparam \macro_inst|controller|serialOutputTrigger[0] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|serialOutputTrigger[0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serialOutputTrigger[0] .BypassEn = 1'b0;
defparam \macro_inst|controller|serialOutputTrigger[0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serialOutputTrigger[1] (
	.A(\macro_inst|controller|serialOutputTrigger [0]),
	.B(\macro_inst|controller|pwmUpdateTrigger~q ),
	.C(vcc),
	.D(\macro_inst|controller|Equal1~2_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serialOutputTrigger [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X51_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serialOutputTrigger[1]~0_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serialOutputTrigger [1]));
defparam \macro_inst|controller|serialOutputTrigger[1] .coord_x = 8;
defparam \macro_inst|controller|serialOutputTrigger[1] .coord_y = 1;
defparam \macro_inst|controller|serialOutputTrigger[1] .coord_z = 3;
defparam \macro_inst|controller|serialOutputTrigger[1] .mask = 16'hF0EC;
defparam \macro_inst|controller|serialOutputTrigger[1] .modeMux = 1'b0;
defparam \macro_inst|controller|serialOutputTrigger[1] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|serialOutputTrigger[1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serialOutputTrigger[1] .BypassEn = 1'b0;
defparam \macro_inst|controller|serialOutputTrigger[1] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serialTrigCounter[0] (
	.A(\macro_inst|controller|Equal1~0_combout ),
	.B(vcc),
	.C(\macro_inst|controller|Equal1~1_combout ),
	.D(\macro_inst|controller|Add0~0_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serialTrigCounter [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X49_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serialTrigCounter~2_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serialTrigCounter [0]));
defparam \macro_inst|controller|serialTrigCounter[0] .coord_x = 6;
defparam \macro_inst|controller|serialTrigCounter[0] .coord_y = 1;
defparam \macro_inst|controller|serialTrigCounter[0] .coord_z = 2;
defparam \macro_inst|controller|serialTrigCounter[0] .mask = 16'h5F00;
defparam \macro_inst|controller|serialTrigCounter[0] .modeMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[0] .BypassEn = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serialTrigCounter[1] (
	.A(vcc),
	.B(\macro_inst|controller|serialTrigCounter [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|Add0~1 ),
	.Qin(\macro_inst|controller|serialTrigCounter [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X49_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|Add0~2_combout ),
	.Cout(\macro_inst|controller|Add0~3 ),
	.Q(\macro_inst|controller|serialTrigCounter [1]));
defparam \macro_inst|controller|serialTrigCounter[1] .coord_x = 6;
defparam \macro_inst|controller|serialTrigCounter[1] .coord_y = 1;
defparam \macro_inst|controller|serialTrigCounter[1] .coord_z = 6;
defparam \macro_inst|controller|serialTrigCounter[1] .mask = 16'h3C3F;
defparam \macro_inst|controller|serialTrigCounter[1] .modeMux = 1'b1;
defparam \macro_inst|controller|serialTrigCounter[1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[1] .BypassEn = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serialTrigCounter[2] (
	.A(\macro_inst|controller|Equal1~0_combout ),
	.B(vcc),
	.C(\macro_inst|controller|Equal1~1_combout ),
	.D(\macro_inst|controller|Add0~4_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serialTrigCounter [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X49_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serialTrigCounter~1_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serialTrigCounter [2]));
defparam \macro_inst|controller|serialTrigCounter[2] .coord_x = 6;
defparam \macro_inst|controller|serialTrigCounter[2] .coord_y = 1;
defparam \macro_inst|controller|serialTrigCounter[2] .coord_z = 13;
defparam \macro_inst|controller|serialTrigCounter[2] .mask = 16'h5F00;
defparam \macro_inst|controller|serialTrigCounter[2] .modeMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[2] .BypassEn = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[2] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serialTrigCounter[3] (
	.A(vcc),
	.B(\macro_inst|controller|serialTrigCounter [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|Add0~5 ),
	.Qin(\macro_inst|controller|serialTrigCounter [3]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X49_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|Add0~6_combout ),
	.Cout(\macro_inst|controller|Add0~7 ),
	.Q(\macro_inst|controller|serialTrigCounter [3]));
defparam \macro_inst|controller|serialTrigCounter[3] .coord_x = 6;
defparam \macro_inst|controller|serialTrigCounter[3] .coord_y = 1;
defparam \macro_inst|controller|serialTrigCounter[3] .coord_z = 8;
defparam \macro_inst|controller|serialTrigCounter[3] .mask = 16'h3C3F;
defparam \macro_inst|controller|serialTrigCounter[3] .modeMux = 1'b1;
defparam \macro_inst|controller|serialTrigCounter[3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[3] .BypassEn = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serialTrigCounter[4] (
	.A(vcc),
	.B(\macro_inst|controller|serialTrigCounter [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|Add0~7 ),
	.Qin(\macro_inst|controller|serialTrigCounter [4]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X49_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|Add0~8_combout ),
	.Cout(\macro_inst|controller|Add0~9 ),
	.Q(\macro_inst|controller|serialTrigCounter [4]));
defparam \macro_inst|controller|serialTrigCounter[4] .coord_x = 6;
defparam \macro_inst|controller|serialTrigCounter[4] .coord_y = 1;
defparam \macro_inst|controller|serialTrigCounter[4] .coord_z = 9;
defparam \macro_inst|controller|serialTrigCounter[4] .mask = 16'hC30C;
defparam \macro_inst|controller|serialTrigCounter[4] .modeMux = 1'b1;
defparam \macro_inst|controller|serialTrigCounter[4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[4] .BypassEn = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serialTrigCounter[5] (
	.A(\macro_inst|controller|Equal1~0_combout ),
	.B(vcc),
	.C(\macro_inst|controller|Add0~10_combout ),
	.D(\macro_inst|controller|Equal1~1_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serialTrigCounter [5]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X49_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serialTrigCounter~0_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serialTrigCounter [5]));
defparam \macro_inst|controller|serialTrigCounter[5] .coord_x = 6;
defparam \macro_inst|controller|serialTrigCounter[5] .coord_y = 1;
defparam \macro_inst|controller|serialTrigCounter[5] .coord_z = 3;
defparam \macro_inst|controller|serialTrigCounter[5] .mask = 16'h50F0;
defparam \macro_inst|controller|serialTrigCounter[5] .modeMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[5] .BypassEn = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serialTrigCounter[6] (
	.A(\macro_inst|controller|serialTrigCounter [6]),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|Add0~11 ),
	.Qin(\macro_inst|controller|serialTrigCounter [6]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X49_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|Add0~12_combout ),
	.Cout(\macro_inst|controller|Add0~13 ),
	.Q(\macro_inst|controller|serialTrigCounter [6]));
defparam \macro_inst|controller|serialTrigCounter[6] .coord_x = 6;
defparam \macro_inst|controller|serialTrigCounter[6] .coord_y = 1;
defparam \macro_inst|controller|serialTrigCounter[6] .coord_z = 11;
defparam \macro_inst|controller|serialTrigCounter[6] .mask = 16'hA50A;
defparam \macro_inst|controller|serialTrigCounter[6] .modeMux = 1'b1;
defparam \macro_inst|controller|serialTrigCounter[6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[6] .BypassEn = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[6] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serialTrigCounter[7] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serialTrigCounter [7]),
	.Cin(\macro_inst|controller|Add0~13 ),
	.Qin(\macro_inst|controller|serialTrigCounter [7]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X49_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|Add0~14_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serialTrigCounter [7]));
defparam \macro_inst|controller|serialTrigCounter[7] .coord_x = 6;
defparam \macro_inst|controller|serialTrigCounter[7] .coord_y = 1;
defparam \macro_inst|controller|serialTrigCounter[7] .coord_z = 12;
defparam \macro_inst|controller|serialTrigCounter[7] .mask = 16'h0FF0;
defparam \macro_inst|controller|serialTrigCounter[7] .modeMux = 1'b1;
defparam \macro_inst|controller|serialTrigCounter[7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[7] .BypassEn = 1'b0;
defparam \macro_inst|controller|serialTrigCounter[7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|Add2~0 (
	.A(\macro_inst|controller|serial|scaler_counter [3]),
	.B(\macro_inst|controller|serial|scaler_counter [1]),
	.C(\macro_inst|controller|serial|scaler_counter [0]),
	.D(\macro_inst|controller|serial|scaler_counter [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|Add2~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|Add2~0 .coord_x = 8;
defparam \macro_inst|controller|serial|Add2~0 .coord_y = 1;
defparam \macro_inst|controller|serial|Add2~0 .coord_z = 0;
defparam \macro_inst|controller|serial|Add2~0 .mask = 16'h6AAA;
defparam \macro_inst|controller|serial|Add2~0 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|Add2~0 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|Add2~0 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|Add2~0 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|Add2~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|Add2~1 (
	.A(vcc),
	.B(\macro_inst|controller|serial|scaler_counter [1]),
	.C(\macro_inst|controller|serial|scaler_counter [0]),
	.D(\macro_inst|controller|serial|scaler_counter [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|Add2~1_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|Add2~1 .coord_x = 8;
defparam \macro_inst|controller|serial|Add2~1 .coord_y = 1;
defparam \macro_inst|controller|serial|Add2~1 .coord_z = 10;
defparam \macro_inst|controller|serial|Add2~1 .mask = 16'h3FC0;
defparam \macro_inst|controller|serial|Add2~1 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|Add2~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|Add2~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|Add2~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|Add2~1 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|Equal0~0 (
	.A(\macro_inst|controller|serial|scaler_counter [3]),
	.B(\macro_inst|controller|serial|scaler_counter [2]),
	.C(\macro_inst|controller|serial|scaler_counter [0]),
	.D(\macro_inst|controller|serial|scaler_counter [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|Equal0~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|Equal0~0 .coord_x = 8;
defparam \macro_inst|controller|serial|Equal0~0 .coord_y = 1;
defparam \macro_inst|controller|serial|Equal0~0 .coord_z = 7;
defparam \macro_inst|controller|serial|Equal0~0 .mask = 16'hFFEF;
defparam \macro_inst|controller|serial|Equal0~0 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|Equal0~0 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|Equal0~0 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|Equal0~0 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|Equal0~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|Equal1~0 (
	.A(\macro_inst|controller|serial|bit_counter [2]),
	.B(\macro_inst|controller|serial|bit_counter [1]),
	.C(\macro_inst|controller|serial|bit_counter [0]),
	.D(\macro_inst|controller|serial|bit_counter [3]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|Equal1~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|Equal1~0 .coord_x = 9;
defparam \macro_inst|controller|serial|Equal1~0 .coord_y = 2;
defparam \macro_inst|controller|serial|Equal1~0 .coord_z = 13;
defparam \macro_inst|controller|serial|Equal1~0 .mask = 16'hFF7F;
defparam \macro_inst|controller|serial|Equal1~0 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|Equal1~0 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|Equal1~0 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|Equal1~0 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|Equal1~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|Equal1~1 (
	.A(\macro_inst|controller|serial|bit_counter [6]),
	.B(\macro_inst|controller|serial|bit_counter [7]),
	.C(\macro_inst|controller|serial|bit_counter [4]),
	.D(\macro_inst|controller|serial|bit_counter [5]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|Equal1~1_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|Equal1~1 .coord_x = 9;
defparam \macro_inst|controller|serial|Equal1~1 .coord_y = 2;
defparam \macro_inst|controller|serial|Equal1~1 .coord_z = 12;
defparam \macro_inst|controller|serial|Equal1~1 .mask = 16'hFFFE;
defparam \macro_inst|controller|serial|Equal1~1 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|Equal1~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|Equal1~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|Equal1~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|Equal1~1 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|Selector2~0 (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.SHIFT~q ),
	.D(\macro_inst|controller|serial|Selector4~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|Selector2~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|Selector2~0 .coord_x = 7;
defparam \macro_inst|controller|serial|Selector2~0 .coord_y = 1;
defparam \macro_inst|controller|serial|Selector2~0 .coord_z = 11;
defparam \macro_inst|controller|serial|Selector2~0 .mask = 16'h00F0;
defparam \macro_inst|controller|serial|Selector2~0 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|Selector2~0 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|Selector2~0 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|Selector2~0 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|Selector2~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|Selector4~0 (
	.A(\macro_inst|controller|serial|byte_counter [1]),
	.B(\macro_inst|controller|serial|byte_counter [0]),
	.C(\macro_inst|controller|serial|byte_counter [3]),
	.D(\macro_inst|controller|serial|byte_counter [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|Selector4~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|Selector4~0 .coord_x = 8;
defparam \macro_inst|controller|serial|Selector4~0 .coord_y = 2;
defparam \macro_inst|controller|serial|Selector4~0 .coord_z = 3;
defparam \macro_inst|controller|serial|Selector4~0 .mask = 16'h0001;
defparam \macro_inst|controller|serial|Selector4~0 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|Selector4~0 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|Selector4~0 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|Selector4~0 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|Selector4~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|Selector4~1 (
	.A(\macro_inst|controller|serial|byte_counter [5]),
	.B(\macro_inst|controller|serial|byte_counter [6]),
	.C(\macro_inst|controller|serial|byte_counter [7]),
	.D(\macro_inst|controller|serial|byte_counter [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|Selector4~1_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|Selector4~1 .coord_x = 8;
defparam \macro_inst|controller|serial|Selector4~1 .coord_y = 2;
defparam \macro_inst|controller|serial|Selector4~1 .coord_z = 14;
defparam \macro_inst|controller|serial|Selector4~1 .mask = 16'h0001;
defparam \macro_inst|controller|serial|Selector4~1 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|Selector4~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|Selector4~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|Selector4~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|Selector4~1 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|Selector4~2 (
	.A(\macro_inst|controller|serial|Equal1~1_combout ),
	.B(\macro_inst|controller|serial|Equal1~0_combout ),
	.C(\macro_inst|controller|serial|Selector4~1_combout ),
	.D(\macro_inst|controller|serial|Selector4~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|Selector4~2_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|Selector4~2 .coord_x = 8;
defparam \macro_inst|controller|serial|Selector4~2 .coord_y = 2;
defparam \macro_inst|controller|serial|Selector4~2 .coord_z = 15;
defparam \macro_inst|controller|serial|Selector4~2 .mask = 16'h1000;
defparam \macro_inst|controller|serial|Selector4~2 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|Selector4~2 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|Selector4~2 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|Selector4~2 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|Selector4~2 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|bit_counter[0] (
	.A(vcc),
	.B(\macro_inst|controller|serial|bit_counter [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|serial|bit_counter [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|bit_counter[7]~8_combout_X50_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|bit_counter[7]~17_combout__SyncReset_X50_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X50_Y2_GND),
	.LutOut(\macro_inst|controller|serial|bit_counter[0]~9_combout ),
	.Cout(\macro_inst|controller|serial|bit_counter[0]~10 ),
	.Q(\macro_inst|controller|serial|bit_counter [0]));
defparam \macro_inst|controller|serial|bit_counter[0] .coord_x = 9;
defparam \macro_inst|controller|serial|bit_counter[0] .coord_y = 2;
defparam \macro_inst|controller|serial|bit_counter[0] .coord_z = 0;
defparam \macro_inst|controller|serial|bit_counter[0] .mask = 16'h33CC;
defparam \macro_inst|controller|serial|bit_counter[0] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[0] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[0] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serial|bit_counter[1] (
	.A(vcc),
	.B(\macro_inst|controller|serial|bit_counter [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|serial|bit_counter[0]~10 ),
	.Qin(\macro_inst|controller|serial|bit_counter [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|bit_counter[7]~8_combout_X50_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|bit_counter[7]~17_combout__SyncReset_X50_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X50_Y2_GND),
	.LutOut(\macro_inst|controller|serial|bit_counter[1]~11_combout ),
	.Cout(\macro_inst|controller|serial|bit_counter[1]~12 ),
	.Q(\macro_inst|controller|serial|bit_counter [1]));
defparam \macro_inst|controller|serial|bit_counter[1] .coord_x = 9;
defparam \macro_inst|controller|serial|bit_counter[1] .coord_y = 2;
defparam \macro_inst|controller|serial|bit_counter[1] .coord_z = 1;
defparam \macro_inst|controller|serial|bit_counter[1] .mask = 16'h3C3F;
defparam \macro_inst|controller|serial|bit_counter[1] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[1] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serial|bit_counter[2] (
	.A(vcc),
	.B(\macro_inst|controller|serial|bit_counter [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|serial|bit_counter[1]~12 ),
	.Qin(\macro_inst|controller|serial|bit_counter [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|bit_counter[7]~8_combout_X50_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|bit_counter[7]~17_combout__SyncReset_X50_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X50_Y2_GND),
	.LutOut(\macro_inst|controller|serial|bit_counter[2]~13_combout ),
	.Cout(\macro_inst|controller|serial|bit_counter[2]~14 ),
	.Q(\macro_inst|controller|serial|bit_counter [2]));
defparam \macro_inst|controller|serial|bit_counter[2] .coord_x = 9;
defparam \macro_inst|controller|serial|bit_counter[2] .coord_y = 2;
defparam \macro_inst|controller|serial|bit_counter[2] .coord_z = 2;
defparam \macro_inst|controller|serial|bit_counter[2] .mask = 16'hC30C;
defparam \macro_inst|controller|serial|bit_counter[2] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[2] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serial|bit_counter[3] (
	.A(vcc),
	.B(\macro_inst|controller|serial|bit_counter [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|serial|bit_counter[2]~14 ),
	.Qin(\macro_inst|controller|serial|bit_counter [3]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|bit_counter[7]~8_combout_X50_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|bit_counter[7]~17_combout__SyncReset_X50_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X50_Y2_GND),
	.LutOut(\macro_inst|controller|serial|bit_counter[3]~15_combout ),
	.Cout(\macro_inst|controller|serial|bit_counter[3]~16 ),
	.Q(\macro_inst|controller|serial|bit_counter [3]));
defparam \macro_inst|controller|serial|bit_counter[3] .coord_x = 9;
defparam \macro_inst|controller|serial|bit_counter[3] .coord_y = 2;
defparam \macro_inst|controller|serial|bit_counter[3] .coord_z = 3;
defparam \macro_inst|controller|serial|bit_counter[3] .mask = 16'h3C3F;
defparam \macro_inst|controller|serial|bit_counter[3] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[3] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serial|bit_counter[4] (
	.A(vcc),
	.B(\macro_inst|controller|serial|bit_counter [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|serial|bit_counter[3]~16 ),
	.Qin(\macro_inst|controller|serial|bit_counter [4]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|bit_counter[7]~8_combout_X50_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|bit_counter[7]~17_combout__SyncReset_X50_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X50_Y2_GND),
	.LutOut(\macro_inst|controller|serial|bit_counter[4]~18_combout ),
	.Cout(\macro_inst|controller|serial|bit_counter[4]~19 ),
	.Q(\macro_inst|controller|serial|bit_counter [4]));
defparam \macro_inst|controller|serial|bit_counter[4] .coord_x = 9;
defparam \macro_inst|controller|serial|bit_counter[4] .coord_y = 2;
defparam \macro_inst|controller|serial|bit_counter[4] .coord_z = 4;
defparam \macro_inst|controller|serial|bit_counter[4] .mask = 16'hC30C;
defparam \macro_inst|controller|serial|bit_counter[4] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[4] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serial|bit_counter[5] (
	.A(vcc),
	.B(\macro_inst|controller|serial|bit_counter [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|serial|bit_counter[4]~19 ),
	.Qin(\macro_inst|controller|serial|bit_counter [5]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|bit_counter[7]~8_combout_X50_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|bit_counter[7]~17_combout__SyncReset_X50_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X50_Y2_GND),
	.LutOut(\macro_inst|controller|serial|bit_counter[5]~20_combout ),
	.Cout(\macro_inst|controller|serial|bit_counter[5]~21 ),
	.Q(\macro_inst|controller|serial|bit_counter [5]));
defparam \macro_inst|controller|serial|bit_counter[5] .coord_x = 9;
defparam \macro_inst|controller|serial|bit_counter[5] .coord_y = 2;
defparam \macro_inst|controller|serial|bit_counter[5] .coord_z = 5;
defparam \macro_inst|controller|serial|bit_counter[5] .mask = 16'h3C3F;
defparam \macro_inst|controller|serial|bit_counter[5] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[5] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[5] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serial|bit_counter[6] (
	.A(vcc),
	.B(\macro_inst|controller|serial|bit_counter [6]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|serial|bit_counter[5]~21 ),
	.Qin(\macro_inst|controller|serial|bit_counter [6]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|bit_counter[7]~8_combout_X50_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|bit_counter[7]~17_combout__SyncReset_X50_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X50_Y2_GND),
	.LutOut(\macro_inst|controller|serial|bit_counter[6]~22_combout ),
	.Cout(\macro_inst|controller|serial|bit_counter[6]~23 ),
	.Q(\macro_inst|controller|serial|bit_counter [6]));
defparam \macro_inst|controller|serial|bit_counter[6] .coord_x = 9;
defparam \macro_inst|controller|serial|bit_counter[6] .coord_y = 2;
defparam \macro_inst|controller|serial|bit_counter[6] .coord_z = 6;
defparam \macro_inst|controller|serial|bit_counter[6] .mask = 16'hC30C;
defparam \macro_inst|controller|serial|bit_counter[6] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[6] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[6] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serial|bit_counter[7] (
	.A(vcc),
	.B(\macro_inst|controller|serial|bit_counter [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|serial|bit_counter[6]~23 ),
	.Qin(\macro_inst|controller|serial|bit_counter [7]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|bit_counter[7]~8_combout_X50_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|bit_counter[7]~17_combout__SyncReset_X50_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X50_Y2_GND),
	.LutOut(\macro_inst|controller|serial|bit_counter[7]~24_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|bit_counter [7]));
defparam \macro_inst|controller|serial|bit_counter[7] .coord_x = 9;
defparam \macro_inst|controller|serial|bit_counter[7] .coord_y = 2;
defparam \macro_inst|controller|serial|bit_counter[7] .coord_z = 7;
defparam \macro_inst|controller|serial|bit_counter[7] .mask = 16'h3C3C;
defparam \macro_inst|controller|serial|bit_counter[7] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[7] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|bit_counter[7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|bit_counter[7]~17 (
	.A(vcc),
	.B(\macro_inst|controller|serial|Equal1~1_combout ),
	.C(\macro_inst|controller|serial|Equal1~0_combout ),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|bit_counter[7]~17_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|bit_counter[7]~17 .coord_x = 8;
defparam \macro_inst|controller|serial|bit_counter[7]~17 .coord_y = 2;
defparam \macro_inst|controller|serial|bit_counter[7]~17 .coord_z = 0;
defparam \macro_inst|controller|serial|bit_counter[7]~17 .mask = 16'h03FF;
defparam \macro_inst|controller|serial|bit_counter[7]~17 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[7]~17 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[7]~17 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[7]~17 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[7]~17 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|bit_counter[7]~8 (
	.A(\macro_inst|controller|serial|state.SHIFT~q ),
	.B(\macro_inst|controller|serial|scaler_counter[0]~0_combout ),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|serial|Equal0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|bit_counter[7]~8_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|bit_counter[7]~8 .coord_x = 8;
defparam \macro_inst|controller|serial|bit_counter[7]~8 .coord_y = 1;
defparam \macro_inst|controller|serial|bit_counter[7]~8 .coord_z = 8;
defparam \macro_inst|controller|serial|bit_counter[7]~8 .mask = 16'h0C8C;
defparam \macro_inst|controller|serial|bit_counter[7]~8 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[7]~8 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[7]~8 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[7]~8 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|bit_counter[7]~8 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|byte_counter[0] (
	.A(vcc),
	.B(\macro_inst|controller|serial|byte_counter [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|serial|byte_counter [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|byte_counter[4]~10_combout_X51_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|state.IDLE~q__SyncReset_X51_Y2_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X51_Y2_GND),
	.LutOut(\macro_inst|controller|serial|byte_counter[0]~8_combout ),
	.Cout(\macro_inst|controller|serial|byte_counter[0]~9 ),
	.Q(\macro_inst|controller|serial|byte_counter [0]));
defparam \macro_inst|controller|serial|byte_counter[0] .coord_x = 8;
defparam \macro_inst|controller|serial|byte_counter[0] .coord_y = 2;
defparam \macro_inst|controller|serial|byte_counter[0] .coord_z = 5;
defparam \macro_inst|controller|serial|byte_counter[0] .mask = 16'h33CC;
defparam \macro_inst|controller|serial|byte_counter[0] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[0] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[0] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serial|byte_counter[1] (
	.A(vcc),
	.B(\macro_inst|controller|serial|byte_counter [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|serial|byte_counter[0]~9 ),
	.Qin(\macro_inst|controller|serial|byte_counter [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|byte_counter[4]~10_combout_X51_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|state.IDLE~q__SyncReset_X51_Y2_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X51_Y2_GND),
	.LutOut(\macro_inst|controller|serial|byte_counter[1]~11_combout ),
	.Cout(\macro_inst|controller|serial|byte_counter[1]~12 ),
	.Q(\macro_inst|controller|serial|byte_counter [1]));
defparam \macro_inst|controller|serial|byte_counter[1] .coord_x = 8;
defparam \macro_inst|controller|serial|byte_counter[1] .coord_y = 2;
defparam \macro_inst|controller|serial|byte_counter[1] .coord_z = 6;
defparam \macro_inst|controller|serial|byte_counter[1] .mask = 16'h3C3F;
defparam \macro_inst|controller|serial|byte_counter[1] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[1] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serial|byte_counter[2] (
	.A(vcc),
	.B(\macro_inst|controller|serial|byte_counter [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|serial|byte_counter[1]~12 ),
	.Qin(\macro_inst|controller|serial|byte_counter [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|byte_counter[4]~10_combout_X51_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|state.IDLE~q__SyncReset_X51_Y2_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X51_Y2_GND),
	.LutOut(\macro_inst|controller|serial|byte_counter[2]~13_combout ),
	.Cout(\macro_inst|controller|serial|byte_counter[2]~14 ),
	.Q(\macro_inst|controller|serial|byte_counter [2]));
defparam \macro_inst|controller|serial|byte_counter[2] .coord_x = 8;
defparam \macro_inst|controller|serial|byte_counter[2] .coord_y = 2;
defparam \macro_inst|controller|serial|byte_counter[2] .coord_z = 7;
defparam \macro_inst|controller|serial|byte_counter[2] .mask = 16'hC30C;
defparam \macro_inst|controller|serial|byte_counter[2] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[2] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serial|byte_counter[3] (
	.A(vcc),
	.B(\macro_inst|controller|serial|byte_counter [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|serial|byte_counter[2]~14 ),
	.Qin(\macro_inst|controller|serial|byte_counter [3]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|byte_counter[4]~10_combout_X51_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|state.IDLE~q__SyncReset_X51_Y2_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X51_Y2_GND),
	.LutOut(\macro_inst|controller|serial|byte_counter[3]~15_combout ),
	.Cout(\macro_inst|controller|serial|byte_counter[3]~16 ),
	.Q(\macro_inst|controller|serial|byte_counter [3]));
defparam \macro_inst|controller|serial|byte_counter[3] .coord_x = 8;
defparam \macro_inst|controller|serial|byte_counter[3] .coord_y = 2;
defparam \macro_inst|controller|serial|byte_counter[3] .coord_z = 8;
defparam \macro_inst|controller|serial|byte_counter[3] .mask = 16'h3C3F;
defparam \macro_inst|controller|serial|byte_counter[3] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[3] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serial|byte_counter[4] (
	.A(vcc),
	.B(\macro_inst|controller|serial|byte_counter [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|serial|byte_counter[3]~16 ),
	.Qin(\macro_inst|controller|serial|byte_counter [4]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|byte_counter[4]~10_combout_X51_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|state.IDLE~q__SyncReset_X51_Y2_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X51_Y2_GND),
	.LutOut(\macro_inst|controller|serial|byte_counter[4]~17_combout ),
	.Cout(\macro_inst|controller|serial|byte_counter[4]~18 ),
	.Q(\macro_inst|controller|serial|byte_counter [4]));
defparam \macro_inst|controller|serial|byte_counter[4] .coord_x = 8;
defparam \macro_inst|controller|serial|byte_counter[4] .coord_y = 2;
defparam \macro_inst|controller|serial|byte_counter[4] .coord_z = 9;
defparam \macro_inst|controller|serial|byte_counter[4] .mask = 16'hC30C;
defparam \macro_inst|controller|serial|byte_counter[4] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[4] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serial|byte_counter[4]~10 (
	.A(\macro_inst|controller|serial|bit_counter[7]~8_combout ),
	.B(\macro_inst|controller|serial|Equal1~1_combout ),
	.C(\macro_inst|controller|serial|Equal1~0_combout ),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|byte_counter[4]~10_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|byte_counter[4]~10 .coord_x = 8;
defparam \macro_inst|controller|serial|byte_counter[4]~10 .coord_y = 2;
defparam \macro_inst|controller|serial|byte_counter[4]~10 .coord_z = 13;
defparam \macro_inst|controller|serial|byte_counter[4]~10 .mask = 16'h02AA;
defparam \macro_inst|controller|serial|byte_counter[4]~10 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[4]~10 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[4]~10 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[4]~10 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[4]~10 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|byte_counter[5] (
	.A(vcc),
	.B(\macro_inst|controller|serial|byte_counter [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|serial|byte_counter[4]~18 ),
	.Qin(\macro_inst|controller|serial|byte_counter [5]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|byte_counter[4]~10_combout_X51_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|state.IDLE~q__SyncReset_X51_Y2_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X51_Y2_GND),
	.LutOut(\macro_inst|controller|serial|byte_counter[5]~19_combout ),
	.Cout(\macro_inst|controller|serial|byte_counter[5]~20 ),
	.Q(\macro_inst|controller|serial|byte_counter [5]));
defparam \macro_inst|controller|serial|byte_counter[5] .coord_x = 8;
defparam \macro_inst|controller|serial|byte_counter[5] .coord_y = 2;
defparam \macro_inst|controller|serial|byte_counter[5] .coord_z = 10;
defparam \macro_inst|controller|serial|byte_counter[5] .mask = 16'h3C3F;
defparam \macro_inst|controller|serial|byte_counter[5] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[5] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[5] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serial|byte_counter[6] (
	.A(vcc),
	.B(\macro_inst|controller|serial|byte_counter [6]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|serial|byte_counter[5]~20 ),
	.Qin(\macro_inst|controller|serial|byte_counter [6]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|byte_counter[4]~10_combout_X51_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|state.IDLE~q__SyncReset_X51_Y2_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X51_Y2_GND),
	.LutOut(\macro_inst|controller|serial|byte_counter[6]~21_combout ),
	.Cout(\macro_inst|controller|serial|byte_counter[6]~22 ),
	.Q(\macro_inst|controller|serial|byte_counter [6]));
defparam \macro_inst|controller|serial|byte_counter[6] .coord_x = 8;
defparam \macro_inst|controller|serial|byte_counter[6] .coord_y = 2;
defparam \macro_inst|controller|serial|byte_counter[6] .coord_z = 11;
defparam \macro_inst|controller|serial|byte_counter[6] .mask = 16'hC30C;
defparam \macro_inst|controller|serial|byte_counter[6] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[6] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[6] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|serial|byte_counter[7] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|byte_counter [7]),
	.Cin(\macro_inst|controller|serial|byte_counter[6]~22 ),
	.Qin(\macro_inst|controller|serial|byte_counter [7]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|byte_counter[4]~10_combout_X51_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y2_SIG ),
	.SyncReset(\macro_inst|controller|serial|state.IDLE~q__SyncReset_X51_Y2_INV ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X51_Y2_GND),
	.LutOut(\macro_inst|controller|serial|byte_counter[7]~23_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|byte_counter [7]));
defparam \macro_inst|controller|serial|byte_counter[7] .coord_x = 8;
defparam \macro_inst|controller|serial|byte_counter[7] .coord_y = 2;
defparam \macro_inst|controller|serial|byte_counter[7] .coord_z = 12;
defparam \macro_inst|controller|serial|byte_counter[7] .mask = 16'h0FF0;
defparam \macro_inst|controller|serial|byte_counter[7] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|byte_counter[7] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|byte_counter[7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|scaler_counter[0] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|serial|scaler_counter [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|scaler_counter[0]~0_combout_X51_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|scaler_counter~4_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|scaler_counter [0]));
defparam \macro_inst|controller|serial|scaler_counter[0] .coord_x = 8;
defparam \macro_inst|controller|serial|scaler_counter[0] .coord_y = 1;
defparam \macro_inst|controller|serial|scaler_counter[0] .coord_z = 14;
defparam \macro_inst|controller|serial|scaler_counter[0] .mask = 16'h0A0A;
defparam \macro_inst|controller|serial|scaler_counter[0] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[0] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|serial|scaler_counter[0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[0] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|scaler_counter[0]~0 (
	.A(vcc),
	.B(\macro_inst|controller|serialOutputTrigger [1]),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|serialOutputTrigger [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|scaler_counter[0]~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|scaler_counter[0]~0 .coord_x = 8;
defparam \macro_inst|controller|serial|scaler_counter[0]~0 .coord_y = 1;
defparam \macro_inst|controller|serial|scaler_counter[0]~0 .coord_z = 5;
defparam \macro_inst|controller|serial|scaler_counter[0]~0 .mask = 16'hFFFC;
defparam \macro_inst|controller|serial|scaler_counter[0]~0 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[0]~0 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[0]~0 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[0]~0 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[0]~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|scaler_counter[1] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(\macro_inst|controller|serial|scaler_counter [0]),
	.C(vcc),
	.D(\macro_inst|controller|serial|Equal0~0_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|scaler_counter [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|scaler_counter[0]~0_combout_X51_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|scaler_counter~3_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|scaler_counter [1]));
defparam \macro_inst|controller|serial|scaler_counter[1] .coord_x = 8;
defparam \macro_inst|controller|serial|scaler_counter[1] .coord_y = 1;
defparam \macro_inst|controller|serial|scaler_counter[1] .coord_z = 15;
defparam \macro_inst|controller|serial|scaler_counter[1] .mask = 16'h2800;
defparam \macro_inst|controller|serial|scaler_counter[1] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[1] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|serial|scaler_counter[1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[1] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[1] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|scaler_counter[2] (
	.A(\macro_inst|controller|serial|Add2~1_combout ),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|serial|Equal0~0_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|scaler_counter [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|scaler_counter[0]~0_combout_X51_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|scaler_counter~2_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|scaler_counter [2]));
defparam \macro_inst|controller|serial|scaler_counter[2] .coord_x = 8;
defparam \macro_inst|controller|serial|scaler_counter[2] .coord_y = 1;
defparam \macro_inst|controller|serial|scaler_counter[2] .coord_z = 9;
defparam \macro_inst|controller|serial|scaler_counter[2] .mask = 16'hA000;
defparam \macro_inst|controller|serial|scaler_counter[2] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[2] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[2] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|scaler_counter[3] (
	.A(\macro_inst|controller|serial|Add2~0_combout ),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|serial|Equal0~0_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|scaler_counter [3]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|scaler_counter[0]~0_combout_X51_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|scaler_counter~1_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|scaler_counter [3]));
defparam \macro_inst|controller|serial|scaler_counter[3] .coord_x = 8;
defparam \macro_inst|controller|serial|scaler_counter[3] .coord_y = 1;
defparam \macro_inst|controller|serial|scaler_counter[3] .coord_z = 4;
defparam \macro_inst|controller|serial|scaler_counter[3] .mask = 16'hA000;
defparam \macro_inst|controller|serial|scaler_counter[3] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[3] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|scaler_counter[3] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data [168]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[0]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [0]));
defparam \macro_inst|controller|serial|sdata_reg[0] .coord_x = 20;
defparam \macro_inst|controller|serial|sdata_reg[0] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[0] .coord_z = 1;
defparam \macro_inst|controller|serial|sdata_reg[0] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|sdata_reg[0] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[0] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[0]~0 (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.LOAD~q ),
	.D(\macro_inst|controller|serial|Equal0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[0]~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|sdata_reg[0]~0 .coord_x = 8;
defparam \macro_inst|controller|serial|sdata_reg[0]~0 .coord_y = 1;
defparam \macro_inst|controller|serial|sdata_reg[0]~0 .coord_z = 12;
defparam \macro_inst|controller|serial|sdata_reg[0]~0 .mask = 16'h00F0;
defparam \macro_inst|controller|serial|sdata_reg[0]~0 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[0]~0 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[0]~0 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[0]~0 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[0]~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[10] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data [178]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [10]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[10]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [10]));
defparam \macro_inst|controller|serial|sdata_reg[10] .coord_x = 20;
defparam \macro_inst|controller|serial|sdata_reg[10] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[10] .coord_z = 11;
defparam \macro_inst|controller|serial|sdata_reg[10] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|sdata_reg[10] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[10] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[10] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[11] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data [179]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [11]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[11]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [11]));
defparam \macro_inst|controller|serial|sdata_reg[11] .coord_x = 11;
defparam \macro_inst|controller|serial|sdata_reg[11] .coord_y = 1;
defparam \macro_inst|controller|serial|sdata_reg[11] .coord_z = 3;
defparam \macro_inst|controller|serial|sdata_reg[11] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|sdata_reg[11] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[11] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[11] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[12] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [180]),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [12]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(SyncReset_X52_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X52_Y2_VCC),
	.LutOut(\~GND~combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [12]));
defparam \macro_inst|controller|serial|sdata_reg[12] .coord_x = 16;
defparam \macro_inst|controller|serial|sdata_reg[12] .coord_y = 5;
defparam \macro_inst|controller|serial|sdata_reg[12] .coord_z = 0;
defparam \macro_inst|controller|serial|sdata_reg[12] .mask = 16'h0000;
defparam \macro_inst|controller|serial|sdata_reg[12] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[12] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|sdata_reg[12] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[13] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data [181]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [13]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[13]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [13]));
defparam \macro_inst|controller|serial|sdata_reg[13] .coord_x = 20;
defparam \macro_inst|controller|serial|sdata_reg[13] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[13] .coord_z = 9;
defparam \macro_inst|controller|serial|sdata_reg[13] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|sdata_reg[13] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[13] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[13] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[14] (
	.A(),
	.B(),
	.C(\macro_inst|controller|serial|shift_data [182]),
	.D(),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [14]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(SyncReset_X51_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X51_Y4_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [14]));
defparam \macro_inst|controller|serial|sdata_reg[14] .coord_x = 15;
defparam \macro_inst|controller|serial|sdata_reg[14] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[14] .coord_z = 10;
defparam \macro_inst|controller|serial|sdata_reg[14] .mask = 16'hFFFF;
defparam \macro_inst|controller|serial|sdata_reg[14] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|sdata_reg[14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[14] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|sdata_reg[14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[15] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data [183]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [15]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[15]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [15]));
defparam \macro_inst|controller|serial|sdata_reg[15] .coord_x = 20;
defparam \macro_inst|controller|serial|sdata_reg[15] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[15] .coord_z = 0;
defparam \macro_inst|controller|serial|sdata_reg[15] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|sdata_reg[15] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[15] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[16] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [184]),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [16]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[16]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [16]));
defparam \macro_inst|controller|serial|sdata_reg[16] .coord_x = 20;
defparam \macro_inst|controller|serial|sdata_reg[16] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[16] .coord_z = 14;
defparam \macro_inst|controller|serial|sdata_reg[16] .mask = 16'hF0F0;
defparam \macro_inst|controller|serial|sdata_reg[16] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[16] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[16] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[16] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[16] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[17] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data [185]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [17]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[17]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [17]));
defparam \macro_inst|controller|serial|sdata_reg[17] .coord_x = 20;
defparam \macro_inst|controller|serial|sdata_reg[17] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[17] .coord_z = 6;
defparam \macro_inst|controller|serial|sdata_reg[17] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|sdata_reg[17] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[17] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[17] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[17] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[17] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[18] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data [186]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [18]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[18]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [18]));
defparam \macro_inst|controller|serial|sdata_reg[18] .coord_x = 20;
defparam \macro_inst|controller|serial|sdata_reg[18] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[18] .coord_z = 5;
defparam \macro_inst|controller|serial|sdata_reg[18] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|sdata_reg[18] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[18] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[18] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[18] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[18] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[19] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [187]),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [19]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[19]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [19]));
defparam \macro_inst|controller|serial|sdata_reg[19] .coord_x = 20;
defparam \macro_inst|controller|serial|sdata_reg[19] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[19] .coord_z = 3;
defparam \macro_inst|controller|serial|sdata_reg[19] .mask = 16'hF0F0;
defparam \macro_inst|controller|serial|sdata_reg[19] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[19] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[19] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[19] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[19] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[1] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data [169]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[1]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [1]));
defparam \macro_inst|controller|serial|sdata_reg[1] .coord_x = 16;
defparam \macro_inst|controller|serial|sdata_reg[1] .coord_y = 5;
defparam \macro_inst|controller|serial|sdata_reg[1] .coord_z = 9;
defparam \macro_inst|controller|serial|sdata_reg[1] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|sdata_reg[1] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[1] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[1] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[20] (
	.A(\macro_inst|controller|serial|shift_data [162]),
	.B(\macro_inst|controller|sm_pwm|data [186]),
	.C(\macro_inst|controller|serial|shift_data [188]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [20]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(SyncReset_X53_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X53_Y4_VCC),
	.LutOut(\macro_inst|controller|serial|shift_data~11_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [20]));
defparam \macro_inst|controller|serial|sdata_reg[20] .coord_x = 15;
defparam \macro_inst|controller|serial|sdata_reg[20] .coord_y = 4;
defparam \macro_inst|controller|serial|sdata_reg[20] .coord_z = 11;
defparam \macro_inst|controller|serial|sdata_reg[20] .mask = 16'hAA33;
defparam \macro_inst|controller|serial|sdata_reg[20] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[20] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[20] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[20] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|sdata_reg[20] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[21] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data [189]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [21]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[21]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [21]));
defparam \macro_inst|controller|serial|sdata_reg[21] .coord_x = 20;
defparam \macro_inst|controller|serial|sdata_reg[21] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[21] .coord_z = 12;
defparam \macro_inst|controller|serial|sdata_reg[21] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|sdata_reg[21] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[21] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[21] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[21] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[21] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[22] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(\macro_inst|controller|serial|shift_data [86]),
	.C(\macro_inst|controller|serial|shift_data [190]),
	.D(\macro_inst|controller|sm_pwm|data [110]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [22]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(SyncReset_X51_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X51_Y4_VCC),
	.LutOut(\macro_inst|controller|serial|shift_data~79_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [22]));
defparam \macro_inst|controller|serial|sdata_reg[22] .coord_x = 15;
defparam \macro_inst|controller|serial|sdata_reg[22] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[22] .coord_z = 12;
defparam \macro_inst|controller|serial|sdata_reg[22] .mask = 16'h88DD;
defparam \macro_inst|controller|serial|sdata_reg[22] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[22] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[22] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[22] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|sdata_reg[22] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[23] (
	.A(),
	.B(),
	.C(\macro_inst|controller|serial|shift_data [191]),
	.D(),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [23]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ),
	.SyncReset(SyncReset_X54_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y1_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [23]));
defparam \macro_inst|controller|serial|sdata_reg[23] .coord_x = 20;
defparam \macro_inst|controller|serial|sdata_reg[23] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[23] .coord_z = 7;
defparam \macro_inst|controller|serial|sdata_reg[23] .mask = 16'hFFFF;
defparam \macro_inst|controller|serial|sdata_reg[23] .modeMux = 1'b1;
defparam \macro_inst|controller|serial|sdata_reg[23] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[23] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[23] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|sdata_reg[23] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[2] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data [170]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[2]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [2]));
defparam \macro_inst|controller|serial|sdata_reg[2] .coord_x = 20;
defparam \macro_inst|controller|serial|sdata_reg[2] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[2] .coord_z = 10;
defparam \macro_inst|controller|serial|sdata_reg[2] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|sdata_reg[2] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[2] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[2] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[3] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data [171]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [3]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[3]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [3]));
defparam \macro_inst|controller|serial|sdata_reg[3] .coord_x = 20;
defparam \macro_inst|controller|serial|sdata_reg[3] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[3] .coord_z = 13;
defparam \macro_inst|controller|serial|sdata_reg[3] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|sdata_reg[3] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[3] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[3] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[4] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(\macro_inst|controller|sm_pwm|data [185]),
	.C(\macro_inst|controller|serial|shift_data [172]),
	.D(\macro_inst|controller|serial|shift_data [161]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [4]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(SyncReset_X53_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X53_Y4_VCC),
	.LutOut(\macro_inst|controller|serial|shift_data~10_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [4]));
defparam \macro_inst|controller|serial|sdata_reg[4] .coord_x = 15;
defparam \macro_inst|controller|serial|sdata_reg[4] .coord_y = 4;
defparam \macro_inst|controller|serial|sdata_reg[4] .coord_z = 13;
defparam \macro_inst|controller|serial|sdata_reg[4] .mask = 16'hBB11;
defparam \macro_inst|controller|serial|sdata_reg[4] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[4] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|sdata_reg[4] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[5] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [173]),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [5]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[5]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [5]));
defparam \macro_inst|controller|serial|sdata_reg[5] .coord_x = 20;
defparam \macro_inst|controller|serial|sdata_reg[5] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[5] .coord_z = 15;
defparam \macro_inst|controller|serial|sdata_reg[5] .mask = 16'hF0F0;
defparam \macro_inst|controller|serial|sdata_reg[5] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[5] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[6] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [174]),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [6]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X54_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[6]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [6]));
defparam \macro_inst|controller|serial|sdata_reg[6] .coord_x = 20;
defparam \macro_inst|controller|serial|sdata_reg[6] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[6] .coord_z = 2;
defparam \macro_inst|controller|serial|sdata_reg[6] .mask = 16'hF0F0;
defparam \macro_inst|controller|serial|sdata_reg[6] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[6] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[7] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data [175]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [7]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[7]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [7]));
defparam \macro_inst|controller|serial|sdata_reg[7] .coord_x = 11;
defparam \macro_inst|controller|serial|sdata_reg[7] .coord_y = 1;
defparam \macro_inst|controller|serial|sdata_reg[7] .coord_z = 4;
defparam \macro_inst|controller|serial|sdata_reg[7] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|sdata_reg[7] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[7] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[8] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data [176]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [8]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[8]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [8]));
defparam \macro_inst|controller|serial|sdata_reg[8] .coord_x = 11;
defparam \macro_inst|controller|serial|sdata_reg[8] .coord_y = 1;
defparam \macro_inst|controller|serial|sdata_reg[8] .coord_z = 14;
defparam \macro_inst|controller|serial|sdata_reg[8] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|sdata_reg[8] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[8] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[8] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sdata_reg[9] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data [177]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sdata_reg [9]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|sdata_reg[0]~0_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sdata_reg[9]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sdata_reg [9]));
defparam \macro_inst|controller|serial|sdata_reg[9] .coord_x = 15;
defparam \macro_inst|controller|serial|sdata_reg[9] .coord_y = 2;
defparam \macro_inst|controller|serial|sdata_reg[9] .coord_z = 0;
defparam \macro_inst|controller|serial|sdata_reg[9] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|sdata_reg[9] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[9] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sdata_reg[9] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shi (
	.A(\macro_inst|controller|serial|state.SHIFT~q ),
	.B(\macro_inst|controller|serial|shi~0_combout ),
	.C(vcc),
	.D(\macro_inst|controller|serial|state.LATCH~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shi~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X50_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shi~1_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shi~q ));
defparam \macro_inst|controller|serial|shi .coord_x = 7;
defparam \macro_inst|controller|serial|shi .coord_y = 1;
defparam \macro_inst|controller|serial|shi .coord_z = 13;
defparam \macro_inst|controller|serial|shi .mask = 16'hF8B8;
defparam \macro_inst|controller|serial|shi .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shi .FeedbackMux = 1'b1;
defparam \macro_inst|controller|serial|shi .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shi .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shi .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[0] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [0]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~169_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [0]));
defparam \macro_inst|controller|serial|shift_data[0] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[0] .coord_y = 9;
defparam \macro_inst|controller|serial|shift_data[0] .coord_z = 0;
defparam \macro_inst|controller|serial|shift_data[0] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[0] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[0] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[100] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [76]),
	.C(\macro_inst|controller|sm_pwm|data [100]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [100]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~91_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [100]));
defparam \macro_inst|controller|serial|shift_data[100] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[100] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[100] .coord_z = 10;
defparam \macro_inst|controller|serial|shift_data[100] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[100] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[100] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[100] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[100] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[100] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[101] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [77]),
	.C(\macro_inst|controller|sm_pwm|data [101]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [101]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~92_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [101]));
defparam \macro_inst|controller|serial|shift_data[101] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[101] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[101] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[101] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[101] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[101] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[101] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[101] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[101] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[102] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [102]),
	.C(\macro_inst|controller|serial|shift_data [78]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [102]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~93_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [102]));
defparam \macro_inst|controller|serial|shift_data[102] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[102] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[102] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[102] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[102] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[102] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[102] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[102] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[102] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[103] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [79]),
	.C(\macro_inst|controller|sm_pwm|data [103]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [103]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~94_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [103]));
defparam \macro_inst|controller|serial|shift_data[103] .coord_x = 18;
defparam \macro_inst|controller|serial|shift_data[103] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[103] .coord_z = 7;
defparam \macro_inst|controller|serial|shift_data[103] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[103] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[103] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[103] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[103] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[103] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[104] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [104]),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|serial|shift_data [80]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [104]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~95_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [104]));
defparam \macro_inst|controller|serial|shift_data[104] .coord_x = 11;
defparam \macro_inst|controller|serial|shift_data[104] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[104] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[104] .mask = 16'hF303;
defparam \macro_inst|controller|serial|shift_data[104] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[104] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[104] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[104] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[104] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[105] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [81]),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [105]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [105]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~96_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [105]));
defparam \macro_inst|controller|serial|shift_data[105] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[105] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[105] .coord_z = 14;
defparam \macro_inst|controller|serial|shift_data[105] .mask = 16'hC0CF;
defparam \macro_inst|controller|serial|shift_data[105] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[105] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[105] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[105] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[105] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[106] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [82]),
	.C(\macro_inst|controller|sm_pwm|data [106]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [106]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~75_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [106]));
defparam \macro_inst|controller|serial|shift_data[106] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[106] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[106] .coord_z = 8;
defparam \macro_inst|controller|serial|shift_data[106] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[106] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[106] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[106] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[106] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[106] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[107] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [83]),
	.C(\macro_inst|controller|sm_pwm|data [107]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [107]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~76_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [107]));
defparam \macro_inst|controller|serial|shift_data[107] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[107] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[107] .coord_z = 13;
defparam \macro_inst|controller|serial|shift_data[107] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[107] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[107] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[107] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[107] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[107] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[108] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [84]),
	.C(\macro_inst|controller|sm_pwm|data [108]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [108]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~77_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [108]));
defparam \macro_inst|controller|serial|shift_data[108] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[108] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[108] .coord_z = 14;
defparam \macro_inst|controller|serial|shift_data[108] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[108] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[108] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[108] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[108] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[108] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[109] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [85]),
	.C(\macro_inst|controller|sm_pwm|data [109]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [109]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~78_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [109]));
defparam \macro_inst|controller|serial|shift_data[109] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[109] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[109] .coord_z = 5;
defparam \macro_inst|controller|serial|shift_data[109] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[109] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[109] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[109] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[109] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[109] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[10] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [10]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [10]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~171_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [10]));
defparam \macro_inst|controller|serial|shift_data[10] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[10] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[10] .coord_z = 1;
defparam \macro_inst|controller|serial|shift_data[10] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[10] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[10] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[10] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[110] (
	.A(\macro_inst|controller|sm_pwm|data [133]),
	.B(\macro_inst|controller|serial|shift_data [109]),
	.C(\macro_inst|controller|serial|shift_data~79_combout ),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [110]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(SyncReset_X52_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X52_Y4_VCC),
	.LutOut(\macro_inst|controller|serial|shift_data~54_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [110]));
defparam \macro_inst|controller|serial|shift_data[110] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[110] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[110] .coord_z = 12;
defparam \macro_inst|controller|serial|shift_data[110] .mask = 16'hCC55;
defparam \macro_inst|controller|serial|shift_data[110] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[110] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[110] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[110] .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|shift_data[110] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[111] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [87]),
	.C(\macro_inst|controller|sm_pwm|data [111]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [111]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~80_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [111]));
defparam \macro_inst|controller|serial|shift_data[111] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[111] .coord_y = 10;
defparam \macro_inst|controller|serial|shift_data[111] .coord_z = 11;
defparam \macro_inst|controller|serial|shift_data[111] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[111] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[111] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[111] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[111] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[111] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[112] (
	.A(\macro_inst|controller|serial|shift_data [88]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [112]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [112]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~81_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [112]));
defparam \macro_inst|controller|serial|shift_data[112] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[112] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[112] .coord_z = 9;
defparam \macro_inst|controller|serial|shift_data[112] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[112] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[112] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[112] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[112] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[112] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[113] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [89]),
	.C(\macro_inst|controller|sm_pwm|data [113]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [113]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~82_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [113]));
defparam \macro_inst|controller|serial|shift_data[113] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[113] .coord_y = 4;
defparam \macro_inst|controller|serial|shift_data[113] .coord_z = 9;
defparam \macro_inst|controller|serial|shift_data[113] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[113] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[113] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[113] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[113] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[113] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[114] (
	.A(\macro_inst|controller|serial|shift_data [90]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [114]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [114]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~83_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [114]));
defparam \macro_inst|controller|serial|shift_data[114] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[114] .coord_y = 4;
defparam \macro_inst|controller|serial|shift_data[114] .coord_z = 14;
defparam \macro_inst|controller|serial|shift_data[114] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[114] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[114] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[114] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[114] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[114] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[115] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [115]),
	.C(\macro_inst|controller|serial|shift_data [91]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [115]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~84_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [115]));
defparam \macro_inst|controller|serial|shift_data[115] .coord_x = 18;
defparam \macro_inst|controller|serial|shift_data[115] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[115] .coord_z = 3;
defparam \macro_inst|controller|serial|shift_data[115] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[115] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[115] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[115] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[115] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[115] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[116] (
	.A(\macro_inst|controller|serial|shift_data [92]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [116]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [116]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~86_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [116]));
defparam \macro_inst|controller|serial|shift_data[116] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[116] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[116] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[116] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[116] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[116] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[116] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[116] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[116] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[117] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [117]),
	.C(\macro_inst|controller|serial|shift_data [93]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [117]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~87_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [117]));
defparam \macro_inst|controller|serial|shift_data[117] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[117] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[117] .coord_z = 8;
defparam \macro_inst|controller|serial|shift_data[117] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[117] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[117] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[117] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[117] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[117] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[118] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [118]),
	.C(\macro_inst|controller|serial|shift_data [94]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [118]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~88_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [118]));
defparam \macro_inst|controller|serial|shift_data[118] .coord_x = 14;
defparam \macro_inst|controller|serial|shift_data[118] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[118] .coord_z = 0;
defparam \macro_inst|controller|serial|shift_data[118] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[118] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[118] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[118] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[118] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[118] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[119] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [95]),
	.C(\macro_inst|controller|sm_pwm|data [119]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [119]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~89_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [119]));
defparam \macro_inst|controller|serial|shift_data[119] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[119] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[119] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[119] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[119] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[119] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[119] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[119] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[119] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[11] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [11]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [11]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~172_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [11]));
defparam \macro_inst|controller|serial|shift_data[11] .coord_x = 11;
defparam \macro_inst|controller|serial|shift_data[11] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[11] .coord_z = 13;
defparam \macro_inst|controller|serial|shift_data[11] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[11] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[11] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[11] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[120] (
	.A(\macro_inst|controller|serial|shift_data [96]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [120]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [120]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~49_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [120]));
defparam \macro_inst|controller|serial|shift_data[120] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[120] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[120] .coord_z = 11;
defparam \macro_inst|controller|serial|shift_data[120] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[120] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[120] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[120] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[120] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[120] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[121] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [121]),
	.C(\macro_inst|controller|serial|shift_data [97]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [121]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~50_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [121]));
defparam \macro_inst|controller|serial|shift_data[121] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[121] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[121] .coord_z = 6;
defparam \macro_inst|controller|serial|shift_data[121] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[121] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[121] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[121] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[121] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[121] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[122] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [122]),
	.C(\macro_inst|controller|serial|shift_data [98]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [122]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~61_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [122]));
defparam \macro_inst|controller|serial|shift_data[122] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[122] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[122] .coord_z = 11;
defparam \macro_inst|controller|serial|shift_data[122] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[122] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[122] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[122] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[122] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[122] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[123] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [99]),
	.C(\macro_inst|controller|sm_pwm|data [123]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [123]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~66_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [123]));
defparam \macro_inst|controller|serial|shift_data[123] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[123] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[123] .coord_z = 11;
defparam \macro_inst|controller|serial|shift_data[123] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[123] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[123] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[123] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[123] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[123] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[124] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [100]),
	.C(\macro_inst|controller|sm_pwm|data [124]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [124]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~67_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [124]));
defparam \macro_inst|controller|serial|shift_data[124] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[124] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[124] .coord_z = 11;
defparam \macro_inst|controller|serial|shift_data[124] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[124] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[124] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[124] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[124] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[124] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[125] (
	.A(\macro_inst|controller|serial|shift_data [101]),
	.B(\macro_inst|controller|serial|state.IDLE~q ),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|data [125]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [125]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~68_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [125]));
defparam \macro_inst|controller|serial|shift_data[125] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[125] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[125] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[125] .mask = 16'h88BB;
defparam \macro_inst|controller|serial|shift_data[125] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[125] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[125] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[125] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[125] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[126] (
	.A(\macro_inst|controller|sm_pwm|data [126]),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [102]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [126]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~69_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [126]));
defparam \macro_inst|controller|serial|shift_data[126] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[126] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[126] .coord_z = 14;
defparam \macro_inst|controller|serial|shift_data[126] .mask = 16'hF055;
defparam \macro_inst|controller|serial|shift_data[126] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[126] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[126] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[126] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[126] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[127] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [103]),
	.C(\macro_inst|controller|sm_pwm|data [127]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [127]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~70_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [127]));
defparam \macro_inst|controller|serial|shift_data[127] .coord_x = 18;
defparam \macro_inst|controller|serial|shift_data[127] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[127] .coord_z = 4;
defparam \macro_inst|controller|serial|shift_data[127] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[127] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[127] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[127] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[127] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[127] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[128] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [104]),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [128]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [128]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~71_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [128]));
defparam \macro_inst|controller|serial|shift_data[128] .coord_x = 11;
defparam \macro_inst|controller|serial|shift_data[128] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[128] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[128] .mask = 16'hC0CF;
defparam \macro_inst|controller|serial|shift_data[128] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[128] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[128] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[128] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[128] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[129] (
	.A(\macro_inst|controller|serial|shift_data [105]),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [129]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [129]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~72_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [129]));
defparam \macro_inst|controller|serial|shift_data[129] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[129] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[129] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[129] .mask = 16'hA0AF;
defparam \macro_inst|controller|serial|shift_data[129] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[129] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[129] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[129] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[129] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[12] (
	.A(\macro_inst|controller|sm_pwm|data [12]),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [12]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~173_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [12]));
defparam \macro_inst|controller|serial|shift_data[12] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[12] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[12] .coord_z = 1;
defparam \macro_inst|controller|serial|shift_data[12] .mask = 16'h0055;
defparam \macro_inst|controller|serial|shift_data[12] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[12] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[12] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[130] (
	.A(\macro_inst|controller|serial|shift_data [106]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [130]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [130]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~51_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [130]));
defparam \macro_inst|controller|serial|shift_data[130] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[130] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[130] .coord_z = 0;
defparam \macro_inst|controller|serial|shift_data[130] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[130] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[130] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[130] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[130] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[130] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[131] (
	.A(\macro_inst|controller|sm_pwm|data [131]),
	.B(\macro_inst|controller|serial|shift_data [107]),
	.C(vcc),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [131]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~52_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [131]));
defparam \macro_inst|controller|serial|shift_data[131] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[131] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[131] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[131] .mask = 16'hCC55;
defparam \macro_inst|controller|serial|shift_data[131] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[131] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[131] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[131] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[131] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[132] (
	.A(\macro_inst|controller|serial|shift_data [108]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [132]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [132]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~53_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [132]));
defparam \macro_inst|controller|serial|shift_data[132] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[132] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[132] .coord_z = 7;
defparam \macro_inst|controller|serial|shift_data[132] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[132] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[132] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[132] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[132] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[132] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[133] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data~54_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [133]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data[133]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [133]));
defparam \macro_inst|controller|serial|shift_data[133] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[133] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[133] .coord_z = 12;
defparam \macro_inst|controller|serial|shift_data[133] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|shift_data[133] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[133] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[133] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[133] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[133] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[134] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [134]),
	.D(\macro_inst|controller|serial|shift_data [110]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [134]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~55_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [134]));
defparam \macro_inst|controller|serial|shift_data[134] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[134] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[134] .coord_z = 6;
defparam \macro_inst|controller|serial|shift_data[134] .mask = 16'hAF05;
defparam \macro_inst|controller|serial|shift_data[134] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[134] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[134] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[134] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[134] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[135] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [111]),
	.C(\macro_inst|controller|sm_pwm|data [135]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [135]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~56_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [135]));
defparam \macro_inst|controller|serial|shift_data[135] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[135] .coord_y = 10;
defparam \macro_inst|controller|serial|shift_data[135] .coord_z = 14;
defparam \macro_inst|controller|serial|shift_data[135] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[135] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[135] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[135] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[135] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[135] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[136] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [112]),
	.C(\macro_inst|controller|sm_pwm|data [136]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [136]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~57_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [136]));
defparam \macro_inst|controller|serial|shift_data[136] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[136] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[136] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[136] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[136] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[136] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[136] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[136] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[136] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[137] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [113]),
	.C(\macro_inst|controller|sm_pwm|data [137]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [137]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~58_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [137]));
defparam \macro_inst|controller|serial|shift_data[137] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[137] .coord_y = 4;
defparam \macro_inst|controller|serial|shift_data[137] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[137] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[137] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[137] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[137] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[137] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[137] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[138] (
	.A(\macro_inst|controller|serial|shift_data [114]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [138]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [138]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~59_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [138]));
defparam \macro_inst|controller|serial|shift_data[138] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[138] .coord_y = 4;
defparam \macro_inst|controller|serial|shift_data[138] .coord_z = 5;
defparam \macro_inst|controller|serial|shift_data[138] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[138] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[138] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[138] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[138] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[138] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[139] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [115]),
	.C(\macro_inst|controller|sm_pwm|data [139]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [139]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~60_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [139]));
defparam \macro_inst|controller|serial|shift_data[139] .coord_x = 18;
defparam \macro_inst|controller|serial|shift_data[139] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[139] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[139] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[139] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[139] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[139] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[139] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[139] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[13] (
	.A(vcc),
	.B(\macro_inst|controller|serial|state.IDLE~q ),
	.C(\macro_inst|controller|sm_pwm|data [13]),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [13]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~174_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [13]));
defparam \macro_inst|controller|serial|shift_data[13] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[13] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[13] .coord_z = 3;
defparam \macro_inst|controller|serial|shift_data[13] .mask = 16'h0303;
defparam \macro_inst|controller|serial|shift_data[13] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[13] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[13] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[140] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [116]),
	.C(\macro_inst|controller|sm_pwm|data [140]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [140]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~62_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [140]));
defparam \macro_inst|controller|serial|shift_data[140] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[140] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[140] .coord_z = 3;
defparam \macro_inst|controller|serial|shift_data[140] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[140] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[140] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[140] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[140] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[140] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[141] (
	.A(\macro_inst|controller|serial|shift_data [117]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [141]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [141]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~63_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [141]));
defparam \macro_inst|controller|serial|shift_data[141] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[141] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[141] .coord_z = 14;
defparam \macro_inst|controller|serial|shift_data[141] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[141] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[141] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[141] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[141] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[141] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[142] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [142]),
	.C(\macro_inst|controller|serial|shift_data [118]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [142]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~64_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [142]));
defparam \macro_inst|controller|serial|shift_data[142] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[142] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[142] .coord_z = 9;
defparam \macro_inst|controller|serial|shift_data[142] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[142] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[142] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[142] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[142] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[142] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[143] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [143]),
	.C(\macro_inst|controller|serial|shift_data [119]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [143]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~65_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [143]));
defparam \macro_inst|controller|serial|shift_data[143] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[143] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[143] .coord_z = 11;
defparam \macro_inst|controller|serial|shift_data[143] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[143] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[143] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[143] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[143] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[143] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[144] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [120]),
	.C(\macro_inst|controller|sm_pwm|data [144]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [144]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~25_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [144]));
defparam \macro_inst|controller|serial|shift_data[144] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[144] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[144] .coord_z = 10;
defparam \macro_inst|controller|serial|shift_data[144] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[144] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[144] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[144] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[144] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[144] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[145] (
	.A(vcc),
	.B(\macro_inst|controller|serial|state.IDLE~q ),
	.C(\macro_inst|controller|serial|shift_data [121]),
	.D(\macro_inst|controller|sm_pwm|data [145]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [145]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~26_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [145]));
defparam \macro_inst|controller|serial|shift_data[145] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[145] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[145] .coord_z = 13;
defparam \macro_inst|controller|serial|shift_data[145] .mask = 16'hC0F3;
defparam \macro_inst|controller|serial|shift_data[145] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[145] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[145] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[145] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[145] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[146] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [122]),
	.C(\macro_inst|controller|sm_pwm|data [146]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [146]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~37_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [146]));
defparam \macro_inst|controller|serial|shift_data[146] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[146] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[146] .coord_z = 0;
defparam \macro_inst|controller|serial|shift_data[146] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[146] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[146] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[146] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[146] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[146] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[147] (
	.A(vcc),
	.B(\macro_inst|controller|serial|state.IDLE~q ),
	.C(\macro_inst|controller|sm_pwm|data [147]),
	.D(\macro_inst|controller|serial|shift_data [123]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [147]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~42_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [147]));
defparam \macro_inst|controller|serial|shift_data[147] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[147] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[147] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[147] .mask = 16'hCF03;
defparam \macro_inst|controller|serial|shift_data[147] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[147] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[147] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[147] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[147] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[148] (
	.A(vcc),
	.B(\macro_inst|controller|serial|state.IDLE~q ),
	.C(\macro_inst|controller|sm_pwm|data [148]),
	.D(\macro_inst|controller|serial|shift_data [124]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [148]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~43_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [148]));
defparam \macro_inst|controller|serial|shift_data[148] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[148] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[148] .coord_z = 13;
defparam \macro_inst|controller|serial|shift_data[148] .mask = 16'hCF03;
defparam \macro_inst|controller|serial|shift_data[148] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[148] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[148] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[148] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[148] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[149] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [125]),
	.C(\macro_inst|controller|sm_pwm|data [149]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [149]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~44_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [149]));
defparam \macro_inst|controller|serial|shift_data[149] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[149] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[149] .coord_z = 13;
defparam \macro_inst|controller|serial|shift_data[149] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[149] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[149] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[149] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[149] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[149] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[14] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [14]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [14]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~175_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [14]));
defparam \macro_inst|controller|serial|shift_data[14] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[14] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[14] .coord_z = 1;
defparam \macro_inst|controller|serial|shift_data[14] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[14] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[14] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[150] (
	.A(\macro_inst|controller|sm_pwm|data [150]),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [126]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [150]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~45_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [150]));
defparam \macro_inst|controller|serial|shift_data[150] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[150] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[150] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[150] .mask = 16'hF055;
defparam \macro_inst|controller|serial|shift_data[150] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[150] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[150] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[150] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[150] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[151] (
	.A(\macro_inst|controller|serial|shift_data [127]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [151]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [151]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~46_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [151]));
defparam \macro_inst|controller|serial|shift_data[151] .coord_x = 18;
defparam \macro_inst|controller|serial|shift_data[151] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[151] .coord_z = 1;
defparam \macro_inst|controller|serial|shift_data[151] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[151] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[151] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[151] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[151] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[151] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[152] (
	.A(\macro_inst|controller|serial|shift_data [128]),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [152]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [152]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~47_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [152]));
defparam \macro_inst|controller|serial|shift_data[152] .coord_x = 11;
defparam \macro_inst|controller|serial|shift_data[152] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[152] .coord_z = 12;
defparam \macro_inst|controller|serial|shift_data[152] .mask = 16'hA0AF;
defparam \macro_inst|controller|serial|shift_data[152] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[152] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[152] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[152] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[152] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[153] (
	.A(vcc),
	.B(\macro_inst|controller|serial|state.IDLE~q ),
	.C(\macro_inst|controller|serial|shift_data [129]),
	.D(\macro_inst|controller|sm_pwm|data [153]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [153]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~48_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [153]));
defparam \macro_inst|controller|serial|shift_data[153] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[153] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[153] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[153] .mask = 16'hC0F3;
defparam \macro_inst|controller|serial|shift_data[153] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[153] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[153] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[153] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[153] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[154] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [154]),
	.C(\macro_inst|controller|serial|shift_data [130]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [154]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~27_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [154]));
defparam \macro_inst|controller|serial|shift_data[154] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[154] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[154] .coord_z = 7;
defparam \macro_inst|controller|serial|shift_data[154] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[154] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[154] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[154] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[154] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[154] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[155] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [155]),
	.C(\macro_inst|controller|serial|shift_data [131]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [155]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~28_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [155]));
defparam \macro_inst|controller|serial|shift_data[155] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[155] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[155] .coord_z = 10;
defparam \macro_inst|controller|serial|shift_data[155] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[155] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[155] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[155] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[155] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[155] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[156] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [132]),
	.C(\macro_inst|controller|sm_pwm|data [156]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [156]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~29_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [156]));
defparam \macro_inst|controller|serial|shift_data[156] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[156] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[156] .coord_z = 5;
defparam \macro_inst|controller|serial|shift_data[156] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[156] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[156] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[156] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[156] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[156] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[157] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [133]),
	.C(\macro_inst|controller|sm_pwm|data [157]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [157]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~30_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [157]));
defparam \macro_inst|controller|serial|shift_data[157] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[157] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[157] .coord_z = 5;
defparam \macro_inst|controller|serial|shift_data[157] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[157] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[157] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[157] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[157] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[157] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[158] (
	.A(\macro_inst|controller|serial|shift_data [134]),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [158]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [158]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~31_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [158]));
defparam \macro_inst|controller|serial|shift_data[158] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[158] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[158] .coord_z = 3;
defparam \macro_inst|controller|serial|shift_data[158] .mask = 16'hA0AF;
defparam \macro_inst|controller|serial|shift_data[158] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[158] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[158] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[158] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[158] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[159] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [159]),
	.C(\macro_inst|controller|serial|shift_data [135]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [159]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~32_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [159]));
defparam \macro_inst|controller|serial|shift_data[159] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[159] .coord_y = 10;
defparam \macro_inst|controller|serial|shift_data[159] .coord_z = 4;
defparam \macro_inst|controller|serial|shift_data[159] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[159] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[159] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[159] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[159] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[159] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[15] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [15]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [15]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~176_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [15]));
defparam \macro_inst|controller|serial|shift_data[15] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[15] .coord_y = 10;
defparam \macro_inst|controller|serial|shift_data[15] .coord_z = 5;
defparam \macro_inst|controller|serial|shift_data[15] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[15] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[15] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[160] (
	.A(\macro_inst|controller|serial|shift_data [136]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [160]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [160]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~33_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [160]));
defparam \macro_inst|controller|serial|shift_data[160] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[160] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[160] .coord_z = 0;
defparam \macro_inst|controller|serial|shift_data[160] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[160] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[160] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[160] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[160] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[160] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[161] (
	.A(\macro_inst|controller|sm_pwm|data [161]),
	.B(\macro_inst|controller|serial|shift_data [137]),
	.C(vcc),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [161]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~34_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [161]));
defparam \macro_inst|controller|serial|shift_data[161] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[161] .coord_y = 4;
defparam \macro_inst|controller|serial|shift_data[161] .coord_z = 3;
defparam \macro_inst|controller|serial|shift_data[161] .mask = 16'hCC55;
defparam \macro_inst|controller|serial|shift_data[161] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[161] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[161] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[161] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[161] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[162] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [138]),
	.C(\macro_inst|controller|sm_pwm|data [162]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [162]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~35_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [162]));
defparam \macro_inst|controller|serial|shift_data[162] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[162] .coord_y = 4;
defparam \macro_inst|controller|serial|shift_data[162] .coord_z = 12;
defparam \macro_inst|controller|serial|shift_data[162] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[162] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[162] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[162] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[162] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[162] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[163] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [139]),
	.C(\macro_inst|controller|sm_pwm|data [163]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [163]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~36_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [163]));
defparam \macro_inst|controller|serial|shift_data[163] .coord_x = 18;
defparam \macro_inst|controller|serial|shift_data[163] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[163] .coord_z = 0;
defparam \macro_inst|controller|serial|shift_data[163] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[163] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[163] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[163] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[163] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[163] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[164] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [140]),
	.C(\macro_inst|controller|sm_pwm|data [164]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [164]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~38_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [164]));
defparam \macro_inst|controller|serial|shift_data[164] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[164] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[164] .coord_z = 10;
defparam \macro_inst|controller|serial|shift_data[164] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[164] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[164] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[164] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[164] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[164] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[165] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [165]),
	.C(\macro_inst|controller|serial|shift_data [141]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [165]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~39_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [165]));
defparam \macro_inst|controller|serial|shift_data[165] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[165] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[165] .coord_z = 12;
defparam \macro_inst|controller|serial|shift_data[165] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[165] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[165] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[165] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[165] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[165] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[166] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [142]),
	.C(\macro_inst|controller|sm_pwm|data [166]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [166]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~40_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [166]));
defparam \macro_inst|controller|serial|shift_data[166] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[166] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[166] .coord_z = 4;
defparam \macro_inst|controller|serial|shift_data[166] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[166] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[166] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[166] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[166] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[166] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[167] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [143]),
	.C(\macro_inst|controller|sm_pwm|data [167]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [167]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~41_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [167]));
defparam \macro_inst|controller|serial|shift_data[167] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[167] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[167] .coord_z = 0;
defparam \macro_inst|controller|serial|shift_data[167] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[167] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[167] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[167] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[167] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[167] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[168] (
	.A(\macro_inst|controller|serial|shift_data [144]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [168]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [168]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~0_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [168]));
defparam \macro_inst|controller|serial|shift_data[168] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[168] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[168] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[168] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[168] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[168] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[168] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[168] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[168] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[169] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [145]),
	.C(\macro_inst|controller|sm_pwm|data [169]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [169]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~2_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [169]));
defparam \macro_inst|controller|serial|shift_data[169] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[169] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[169] .coord_z = 3;
defparam \macro_inst|controller|serial|shift_data[169] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[169] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[169] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[169] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[169] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[169] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[16] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [16]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [16]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~177_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [16]));
defparam \macro_inst|controller|serial|shift_data[16] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[16] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[16] .coord_z = 0;
defparam \macro_inst|controller|serial|shift_data[16] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[16] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[16] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[16] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[16] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[16] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[170] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [146]),
	.C(\macro_inst|controller|sm_pwm|data [170]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [170]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~13_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [170]));
defparam \macro_inst|controller|serial|shift_data[170] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[170] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[170] .coord_z = 1;
defparam \macro_inst|controller|serial|shift_data[170] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[170] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[170] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[170] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[170] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[170] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[171] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [171]),
	.C(\macro_inst|controller|serial|shift_data [147]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [171]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~18_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [171]));
defparam \macro_inst|controller|serial|shift_data[171] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[171] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[171] .coord_z = 3;
defparam \macro_inst|controller|serial|shift_data[171] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[171] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[171] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[171] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[171] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[171] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[172] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [172]),
	.C(\macro_inst|controller|serial|shift_data [148]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [172]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~19_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [172]));
defparam \macro_inst|controller|serial|shift_data[172] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[172] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[172] .coord_z = 4;
defparam \macro_inst|controller|serial|shift_data[172] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[172] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[172] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[172] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[172] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[172] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[173] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [149]),
	.C(\macro_inst|controller|sm_pwm|data [173]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [173]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~20_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [173]));
defparam \macro_inst|controller|serial|shift_data[173] .coord_x = 18;
defparam \macro_inst|controller|serial|shift_data[173] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[173] .coord_z = 5;
defparam \macro_inst|controller|serial|shift_data[173] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[173] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[173] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[173] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[173] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[173] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[174] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [150]),
	.C(\macro_inst|controller|sm_pwm|data [174]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [174]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~21_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [174]));
defparam \macro_inst|controller|serial|shift_data[174] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[174] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[174] .coord_z = 4;
defparam \macro_inst|controller|serial|shift_data[174] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[174] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[174] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[174] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[174] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[174] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[175] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [151]),
	.C(\macro_inst|controller|sm_pwm|data [175]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [175]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~22_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [175]));
defparam \macro_inst|controller|serial|shift_data[175] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[175] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[175] .coord_z = 10;
defparam \macro_inst|controller|serial|shift_data[175] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[175] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[175] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[175] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[175] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[175] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[176] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [152]),
	.D(\macro_inst|controller|sm_pwm|data [176]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [176]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~23_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [176]));
defparam \macro_inst|controller|serial|shift_data[176] .coord_x = 11;
defparam \macro_inst|controller|serial|shift_data[176] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[176] .coord_z = 11;
defparam \macro_inst|controller|serial|shift_data[176] .mask = 16'hA0F5;
defparam \macro_inst|controller|serial|shift_data[176] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[176] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[176] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[176] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[176] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[177] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [153]),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [177]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [177]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~24_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [177]));
defparam \macro_inst|controller|serial|shift_data[177] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[177] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[177] .coord_z = 7;
defparam \macro_inst|controller|serial|shift_data[177] .mask = 16'hC0CF;
defparam \macro_inst|controller|serial|shift_data[177] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[177] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[177] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[177] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[177] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[178] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [154]),
	.C(\macro_inst|controller|sm_pwm|data [178]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [178]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~3_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [178]));
defparam \macro_inst|controller|serial|shift_data[178] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[178] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[178] .coord_z = 6;
defparam \macro_inst|controller|serial|shift_data[178] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[178] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[178] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[178] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[178] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[178] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[179] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [179]),
	.C(\macro_inst|controller|serial|shift_data [155]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [179]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~4_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [179]));
defparam \macro_inst|controller|serial|shift_data[179] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[179] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[179] .coord_z = 0;
defparam \macro_inst|controller|serial|shift_data[179] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[179] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[179] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[179] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[179] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[179] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[17] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [17]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [17]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~178_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [17]));
defparam \macro_inst|controller|serial|shift_data[17] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[17] .coord_y = 4;
defparam \macro_inst|controller|serial|shift_data[17] .coord_z = 4;
defparam \macro_inst|controller|serial|shift_data[17] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[17] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[17] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[17] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[17] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[17] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[180] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [156]),
	.C(\macro_inst|controller|sm_pwm|data [180]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [180]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~5_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [180]));
defparam \macro_inst|controller|serial|shift_data[180] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[180] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[180] .coord_z = 4;
defparam \macro_inst|controller|serial|shift_data[180] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[180] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[180] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[180] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[180] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[180] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[181] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [157]),
	.C(\macro_inst|controller|sm_pwm|data [181]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [181]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~6_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [181]));
defparam \macro_inst|controller|serial|shift_data[181] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[181] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[181] .coord_z = 4;
defparam \macro_inst|controller|serial|shift_data[181] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[181] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[181] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[181] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[181] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[181] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[182] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [158]),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [182]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [182]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~7_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [182]));
defparam \macro_inst|controller|serial|shift_data[182] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[182] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[182] .coord_z = 11;
defparam \macro_inst|controller|serial|shift_data[182] .mask = 16'hC0CF;
defparam \macro_inst|controller|serial|shift_data[182] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[182] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[182] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[182] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[182] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[183] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [183]),
	.C(\macro_inst|controller|serial|shift_data [159]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [183]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~8_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [183]));
defparam \macro_inst|controller|serial|shift_data[183] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[183] .coord_y = 10;
defparam \macro_inst|controller|serial|shift_data[183] .coord_z = 8;
defparam \macro_inst|controller|serial|shift_data[183] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[183] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[183] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[183] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[183] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[183] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[184] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [160]),
	.C(\macro_inst|controller|sm_pwm|data [184]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [184]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~9_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [184]));
defparam \macro_inst|controller|serial|shift_data[184] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[184] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[184] .coord_z = 1;
defparam \macro_inst|controller|serial|shift_data[184] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[184] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[184] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[184] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[184] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[184] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[185] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data~10_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [185]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data[185]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [185]));
defparam \macro_inst|controller|serial|shift_data[185] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[185] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[185] .coord_z = 6;
defparam \macro_inst|controller|serial|shift_data[185] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|shift_data[185] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[185] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[185] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[185] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[185] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[186] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|shift_data~11_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [186]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data[186]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [186]));
defparam \macro_inst|controller|serial|shift_data[186] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[186] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[186] .coord_z = 5;
defparam \macro_inst|controller|serial|shift_data[186] .mask = 16'hFF00;
defparam \macro_inst|controller|serial|shift_data[186] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[186] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[186] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[186] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[186] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[187] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [187]),
	.C(\macro_inst|controller|serial|shift_data [163]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [187]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [187]));
defparam \macro_inst|controller|serial|shift_data[187] .coord_x = 18;
defparam \macro_inst|controller|serial|shift_data[187] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[187] .coord_z = 6;
defparam \macro_inst|controller|serial|shift_data[187] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[187] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[187] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[187] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[187] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[187] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[188] (
	.A(\macro_inst|controller|serial|shift_data [164]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [188]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [188]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~14_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [188]));
defparam \macro_inst|controller|serial|shift_data[188] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[188] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[188] .coord_z = 9;
defparam \macro_inst|controller|serial|shift_data[188] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[188] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[188] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[188] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[188] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[188] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[189] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [189]),
	.C(\macro_inst|controller|serial|shift_data [165]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [189]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~15_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [189]));
defparam \macro_inst|controller|serial|shift_data[189] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[189] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[189] .coord_z = 5;
defparam \macro_inst|controller|serial|shift_data[189] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[189] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[189] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[189] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[189] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[189] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[18] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [18]),
	.C(vcc),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [18]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~179_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [18]));
defparam \macro_inst|controller|serial|shift_data[18] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[18] .coord_y = 4;
defparam \macro_inst|controller|serial|shift_data[18] .coord_z = 1;
defparam \macro_inst|controller|serial|shift_data[18] .mask = 16'h0033;
defparam \macro_inst|controller|serial|shift_data[18] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[18] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[18] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[18] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[18] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[190] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [166]),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [190]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [190]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~16_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [190]));
defparam \macro_inst|controller|serial|shift_data[190] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[190] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[190] .coord_z = 13;
defparam \macro_inst|controller|serial|shift_data[190] .mask = 16'hC0CF;
defparam \macro_inst|controller|serial|shift_data[190] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[190] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[190] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[190] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[190] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[191] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [167]),
	.C(\macro_inst|controller|sm_pwm|data [191]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [191]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~17_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [191]));
defparam \macro_inst|controller|serial|shift_data[191] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[191] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[191] .coord_z = 1;
defparam \macro_inst|controller|serial|shift_data[191] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[191] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[191] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[191] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[191] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[191] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[19] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [19]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [19]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~180_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [19]));
defparam \macro_inst|controller|serial|shift_data[19] .coord_x = 17;
defparam \macro_inst|controller|serial|shift_data[19] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[19] .coord_z = 11;
defparam \macro_inst|controller|serial|shift_data[19] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[19] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[19] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[19] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[19] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[19] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[1] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [1]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~170_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [1]));
defparam \macro_inst|controller|serial|shift_data[1] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[1] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[1] .coord_z = 5;
defparam \macro_inst|controller|serial|shift_data[1] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[1] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[1] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[1] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[20] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [20]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [20]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~182_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [20]));
defparam \macro_inst|controller|serial|shift_data[20] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[20] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[20] .coord_z = 13;
defparam \macro_inst|controller|serial|shift_data[20] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[20] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[20] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[20] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[20] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[20] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[21] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [21]),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [21]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~183_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [21]));
defparam \macro_inst|controller|serial|shift_data[21] .coord_x = 14;
defparam \macro_inst|controller|serial|shift_data[21] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[21] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[21] .mask = 16'h0303;
defparam \macro_inst|controller|serial|shift_data[21] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[21] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[21] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[21] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[21] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[22] (
	.A(\macro_inst|controller|sm_pwm|data [22]),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [22]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~184_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [22]));
defparam \macro_inst|controller|serial|shift_data[22] .coord_x = 14;
defparam \macro_inst|controller|serial|shift_data[22] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[22] .coord_z = 3;
defparam \macro_inst|controller|serial|shift_data[22] .mask = 16'h0505;
defparam \macro_inst|controller|serial|shift_data[22] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[22] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[22] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[22] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[22] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[23] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [23]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [23]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~185_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [23]));
defparam \macro_inst|controller|serial|shift_data[23] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[23] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[23] .coord_z = 3;
defparam \macro_inst|controller|serial|shift_data[23] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[23] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[23] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[23] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[23] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[23] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[24] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [0]),
	.D(\macro_inst|controller|sm_pwm|data [24]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [24]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~145_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [24]));
defparam \macro_inst|controller|serial|shift_data[24] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[24] .coord_y = 9;
defparam \macro_inst|controller|serial|shift_data[24] .coord_z = 12;
defparam \macro_inst|controller|serial|shift_data[24] .mask = 16'hA0F5;
defparam \macro_inst|controller|serial|shift_data[24] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[24] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[24] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[24] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[24] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[25] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [1]),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [25]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [25]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~146_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [25]));
defparam \macro_inst|controller|serial|shift_data[25] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[25] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[25] .coord_z = 8;
defparam \macro_inst|controller|serial|shift_data[25] .mask = 16'hC0CF;
defparam \macro_inst|controller|serial|shift_data[25] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[25] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[25] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[25] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[25] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[26] (
	.A(\macro_inst|controller|serial|shift_data [2]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [26]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [26]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~157_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [26]));
defparam \macro_inst|controller|serial|shift_data[26] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[26] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[26] .coord_z = 12;
defparam \macro_inst|controller|serial|shift_data[26] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[26] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[26] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[26] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[26] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[26] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[27] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [3]),
	.C(\macro_inst|controller|sm_pwm|data [27]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [27]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~162_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [27]));
defparam \macro_inst|controller|serial|shift_data[27] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[27] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[27] .coord_z = 7;
defparam \macro_inst|controller|serial|shift_data[27] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[27] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[27] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[27] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[27] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[27] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[28] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [4]),
	.C(\macro_inst|controller|sm_pwm|data [28]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [28]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~163_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [28]));
defparam \macro_inst|controller|serial|shift_data[28] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[28] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[28] .coord_z = 7;
defparam \macro_inst|controller|serial|shift_data[28] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[28] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[28] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[28] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[28] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[28] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[29] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [29]),
	.D(\macro_inst|controller|serial|shift_data [5]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [29]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~164_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [29]));
defparam \macro_inst|controller|serial|shift_data[29] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[29] .coord_y = 9;
defparam \macro_inst|controller|serial|shift_data[29] .coord_z = 3;
defparam \macro_inst|controller|serial|shift_data[29] .mask = 16'hAF05;
defparam \macro_inst|controller|serial|shift_data[29] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[29] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[29] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[29] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[29] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[2] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [2]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~181_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [2]));
defparam \macro_inst|controller|serial|shift_data[2] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[2] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[2] .coord_z = 4;
defparam \macro_inst|controller|serial|shift_data[2] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[2] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[2] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[2] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[30] (
	.A(\macro_inst|controller|sm_pwm|data [30]),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [6]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [30]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~165_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [30]));
defparam \macro_inst|controller|serial|shift_data[30] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[30] .coord_y = 10;
defparam \macro_inst|controller|serial|shift_data[30] .coord_z = 3;
defparam \macro_inst|controller|serial|shift_data[30] .mask = 16'hF055;
defparam \macro_inst|controller|serial|shift_data[30] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[30] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[30] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[30] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[30] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[31] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [7]),
	.C(\macro_inst|controller|sm_pwm|data [31]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [31]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~166_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [31]));
defparam \macro_inst|controller|serial|shift_data[31] .coord_x = 17;
defparam \macro_inst|controller|serial|shift_data[31] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[31] .coord_z = 14;
defparam \macro_inst|controller|serial|shift_data[31] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[31] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[31] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[31] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[31] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[31] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[32] (
	.A(\macro_inst|controller|serial|shift_data [8]),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [32]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [32]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~167_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [32]));
defparam \macro_inst|controller|serial|shift_data[32] .coord_x = 11;
defparam \macro_inst|controller|serial|shift_data[32] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[32] .coord_z = 10;
defparam \macro_inst|controller|serial|shift_data[32] .mask = 16'hA0AF;
defparam \macro_inst|controller|serial|shift_data[32] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[32] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[32] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[32] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[32] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[33] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [9]),
	.C(\macro_inst|controller|sm_pwm|data [33]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [33]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X50_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~168_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [33]));
defparam \macro_inst|controller|serial|shift_data[33] .coord_x = 9;
defparam \macro_inst|controller|serial|shift_data[33] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[33] .coord_z = 7;
defparam \macro_inst|controller|serial|shift_data[33] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[33] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[33] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[33] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[33] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[33] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[34] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [10]),
	.C(\macro_inst|controller|sm_pwm|data [34]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [34]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~147_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [34]));
defparam \macro_inst|controller|serial|shift_data[34] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[34] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[34] .coord_z = 12;
defparam \macro_inst|controller|serial|shift_data[34] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[34] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[34] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[34] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[34] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[34] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[35] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [11]),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [35]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [35]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~148_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [35]));
defparam \macro_inst|controller|serial|shift_data[35] .coord_x = 11;
defparam \macro_inst|controller|serial|shift_data[35] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[35] .coord_z = 9;
defparam \macro_inst|controller|serial|shift_data[35] .mask = 16'hC0CF;
defparam \macro_inst|controller|serial|shift_data[35] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[35] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[35] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[35] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[35] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[36] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [12]),
	.C(\macro_inst|controller|sm_pwm|data [36]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [36]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~149_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [36]));
defparam \macro_inst|controller|serial|shift_data[36] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[36] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[36] .coord_z = 8;
defparam \macro_inst|controller|serial|shift_data[36] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[36] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[36] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[36] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[36] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[36] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[37] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [13]),
	.C(\macro_inst|controller|sm_pwm|data [37]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [37]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~150_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [37]));
defparam \macro_inst|controller|serial|shift_data[37] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[37] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[37] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[37] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[37] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[37] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[37] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[37] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[37] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[38] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [14]),
	.C(\macro_inst|controller|sm_pwm|data [38]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [38]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~151_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [38]));
defparam \macro_inst|controller|serial|shift_data[38] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[38] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[38] .coord_z = 6;
defparam \macro_inst|controller|serial|shift_data[38] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[38] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[38] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[38] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[38] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[38] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[39] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [15]),
	.C(\macro_inst|controller|sm_pwm|data [39]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [39]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~152_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [39]));
defparam \macro_inst|controller|serial|shift_data[39] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[39] .coord_y = 10;
defparam \macro_inst|controller|serial|shift_data[39] .coord_z = 1;
defparam \macro_inst|controller|serial|shift_data[39] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[39] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[39] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[39] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[39] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[39] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[3] (
	.A(\macro_inst|controller|sm_pwm|data [3]),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [3]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~186_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [3]));
defparam \macro_inst|controller|serial|shift_data[3] .coord_x = 11;
defparam \macro_inst|controller|serial|shift_data[3] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[3] .coord_z = 7;
defparam \macro_inst|controller|serial|shift_data[3] .mask = 16'h0505;
defparam \macro_inst|controller|serial|shift_data[3] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[3] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[3] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[40] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [40]),
	.C(\macro_inst|controller|serial|shift_data [16]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [40]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~153_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [40]));
defparam \macro_inst|controller|serial|shift_data[40] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[40] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[40] .coord_z = 1;
defparam \macro_inst|controller|serial|shift_data[40] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[40] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[40] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[40] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[40] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[40] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[41] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [41]),
	.C(\macro_inst|controller|serial|shift_data [17]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [41]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~154_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [41]));
defparam \macro_inst|controller|serial|shift_data[41] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[41] .coord_y = 4;
defparam \macro_inst|controller|serial|shift_data[41] .coord_z = 7;
defparam \macro_inst|controller|serial|shift_data[41] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[41] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[41] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[41] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[41] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[41] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[42] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [18]),
	.C(\macro_inst|controller|sm_pwm|data [42]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [42]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~155_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [42]));
defparam \macro_inst|controller|serial|shift_data[42] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[42] .coord_y = 4;
defparam \macro_inst|controller|serial|shift_data[42] .coord_z = 0;
defparam \macro_inst|controller|serial|shift_data[42] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[42] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[42] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[42] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[42] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[42] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[43] (
	.A(\macro_inst|controller|sm_pwm|data [43]),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [19]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [43]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~156_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [43]));
defparam \macro_inst|controller|serial|shift_data[43] .coord_x = 17;
defparam \macro_inst|controller|serial|shift_data[43] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[43] .coord_z = 10;
defparam \macro_inst|controller|serial|shift_data[43] .mask = 16'hF055;
defparam \macro_inst|controller|serial|shift_data[43] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[43] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[43] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[43] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[43] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[44] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [44]),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|serial|shift_data [20]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [44]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~158_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [44]));
defparam \macro_inst|controller|serial|shift_data[44] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[44] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[44] .coord_z = 8;
defparam \macro_inst|controller|serial|shift_data[44] .mask = 16'hF303;
defparam \macro_inst|controller|serial|shift_data[44] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[44] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[44] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[44] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[44] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[45] (
	.A(\macro_inst|controller|sm_pwm|data [45]),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [21]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [45]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~159_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [45]));
defparam \macro_inst|controller|serial|shift_data[45] .coord_x = 14;
defparam \macro_inst|controller|serial|shift_data[45] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[45] .coord_z = 14;
defparam \macro_inst|controller|serial|shift_data[45] .mask = 16'hF055;
defparam \macro_inst|controller|serial|shift_data[45] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[45] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[45] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[45] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[45] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[46] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [22]),
	.C(\macro_inst|controller|sm_pwm|data [46]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [46]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~160_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [46]));
defparam \macro_inst|controller|serial|shift_data[46] .coord_x = 14;
defparam \macro_inst|controller|serial|shift_data[46] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[46] .coord_z = 1;
defparam \macro_inst|controller|serial|shift_data[46] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[46] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[46] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[46] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[46] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[46] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[47] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [23]),
	.C(\macro_inst|controller|sm_pwm|data [47]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [47]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~161_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [47]));
defparam \macro_inst|controller|serial|shift_data[47] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[47] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[47] .coord_z = 8;
defparam \macro_inst|controller|serial|shift_data[47] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[47] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[47] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[47] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[47] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[47] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[47]~1 (
	.A(\macro_inst|controller|serial|state.LOAD~q ),
	.B(\macro_inst|controller|serial|scaler_counter[0]~0_combout ),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|serial|Equal0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data[47]~1_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|shift_data[47]~1 .coord_x = 8;
defparam \macro_inst|controller|serial|shift_data[47]~1 .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[47]~1 .coord_z = 6;
defparam \macro_inst|controller|serial|shift_data[47]~1 .mask = 16'h0C8C;
defparam \macro_inst|controller|serial|shift_data[47]~1 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[47]~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[47]~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[47]~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[47]~1 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[48] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [24]),
	.D(\macro_inst|controller|sm_pwm|data [48]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [48]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~121_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [48]));
defparam \macro_inst|controller|serial|shift_data[48] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[48] .coord_y = 9;
defparam \macro_inst|controller|serial|shift_data[48] .coord_z = 13;
defparam \macro_inst|controller|serial|shift_data[48] .mask = 16'hA0F5;
defparam \macro_inst|controller|serial|shift_data[48] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[48] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[48] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[48] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[48] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[49] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [25]),
	.C(\macro_inst|controller|sm_pwm|data [49]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [49]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~122_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [49]));
defparam \macro_inst|controller|serial|shift_data[49] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[49] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[49] .coord_z = 8;
defparam \macro_inst|controller|serial|shift_data[49] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[49] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[49] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[49] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[49] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[49] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[4] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [4]),
	.C(vcc),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [4]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~187_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [4]));
defparam \macro_inst|controller|serial|shift_data[4] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[4] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[4] .coord_z = 3;
defparam \macro_inst|controller|serial|shift_data[4] .mask = 16'h0033;
defparam \macro_inst|controller|serial|shift_data[4] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[4] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[4] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[50] (
	.A(\macro_inst|controller|serial|shift_data [26]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [50]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [50]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~133_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [50]));
defparam \macro_inst|controller|serial|shift_data[50] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[50] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[50] .coord_z = 5;
defparam \macro_inst|controller|serial|shift_data[50] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[50] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[50] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[50] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[50] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[50] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[51] (
	.A(\macro_inst|controller|sm_pwm|data [51]),
	.B(\macro_inst|controller|serial|shift_data [27]),
	.C(vcc),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [51]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~138_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [51]));
defparam \macro_inst|controller|serial|shift_data[51] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[51] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[51] .coord_z = 12;
defparam \macro_inst|controller|serial|shift_data[51] .mask = 16'hCC55;
defparam \macro_inst|controller|serial|shift_data[51] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[51] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[51] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[51] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[51] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[52] (
	.A(\macro_inst|controller|sm_pwm|data [52]),
	.B(\macro_inst|controller|serial|shift_data [28]),
	.C(vcc),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [52]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~139_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [52]));
defparam \macro_inst|controller|serial|shift_data[52] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[52] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[52] .coord_z = 9;
defparam \macro_inst|controller|serial|shift_data[52] .mask = 16'hCC55;
defparam \macro_inst|controller|serial|shift_data[52] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[52] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[52] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[52] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[52] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[53] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [29]),
	.D(\macro_inst|controller|sm_pwm|data [53]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [53]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~140_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [53]));
defparam \macro_inst|controller|serial|shift_data[53] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[53] .coord_y = 9;
defparam \macro_inst|controller|serial|shift_data[53] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[53] .mask = 16'hA0F5;
defparam \macro_inst|controller|serial|shift_data[53] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[53] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[53] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[53] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[53] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[54] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [30]),
	.C(\macro_inst|controller|sm_pwm|data [54]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [54]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~141_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [54]));
defparam \macro_inst|controller|serial|shift_data[54] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[54] .coord_y = 10;
defparam \macro_inst|controller|serial|shift_data[54] .coord_z = 10;
defparam \macro_inst|controller|serial|shift_data[54] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[54] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[54] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[54] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[54] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[54] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[55] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [55]),
	.C(\macro_inst|controller|serial|shift_data [31]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [55]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~142_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [55]));
defparam \macro_inst|controller|serial|shift_data[55] .coord_x = 17;
defparam \macro_inst|controller|serial|shift_data[55] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[55] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[55] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[55] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[55] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[55] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[55] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[55] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[56] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [32]),
	.D(\macro_inst|controller|sm_pwm|data [56]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [56]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~143_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [56]));
defparam \macro_inst|controller|serial|shift_data[56] .coord_x = 11;
defparam \macro_inst|controller|serial|shift_data[56] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[56] .coord_z = 5;
defparam \macro_inst|controller|serial|shift_data[56] .mask = 16'hA0F5;
defparam \macro_inst|controller|serial|shift_data[56] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[56] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[56] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[56] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[56] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[57] (
	.A(vcc),
	.B(\macro_inst|controller|serial|state.IDLE~q ),
	.C(\macro_inst|controller|sm_pwm|data [57]),
	.D(\macro_inst|controller|serial|shift_data [33]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [57]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~144_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [57]));
defparam \macro_inst|controller|serial|shift_data[57] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[57] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[57] .coord_z = 4;
defparam \macro_inst|controller|serial|shift_data[57] .mask = 16'hCF03;
defparam \macro_inst|controller|serial|shift_data[57] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[57] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[57] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[57] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[57] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[58] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [34]),
	.C(\macro_inst|controller|sm_pwm|data [58]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [58]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~123_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [58]));
defparam \macro_inst|controller|serial|shift_data[58] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[58] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[58] .coord_z = 13;
defparam \macro_inst|controller|serial|shift_data[58] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[58] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[58] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[58] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[58] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[58] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[59] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [59]),
	.D(\macro_inst|controller|serial|shift_data [35]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [59]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~124_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [59]));
defparam \macro_inst|controller|serial|shift_data[59] .coord_x = 11;
defparam \macro_inst|controller|serial|shift_data[59] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[59] .coord_z = 6;
defparam \macro_inst|controller|serial|shift_data[59] .mask = 16'hAF05;
defparam \macro_inst|controller|serial|shift_data[59] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[59] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[59] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[59] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[59] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[5] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [5]),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [5]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~188_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [5]));
defparam \macro_inst|controller|serial|shift_data[5] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[5] .coord_y = 9;
defparam \macro_inst|controller|serial|shift_data[5] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[5] .mask = 16'h0303;
defparam \macro_inst|controller|serial|shift_data[5] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[5] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[60] (
	.A(\macro_inst|controller|serial|shift_data [36]),
	.B(\macro_inst|controller|serial|state.IDLE~q ),
	.C(\macro_inst|controller|sm_pwm|data [60]),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [60]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~125_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [60]));
defparam \macro_inst|controller|serial|shift_data[60] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[60] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[60] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[60] .mask = 16'h8B8B;
defparam \macro_inst|controller|serial|shift_data[60] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[60] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[60] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[60] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[60] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[61] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [37]),
	.C(\macro_inst|controller|sm_pwm|data [61]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [61]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~126_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [61]));
defparam \macro_inst|controller|serial|shift_data[61] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[61] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[61] .coord_z = 14;
defparam \macro_inst|controller|serial|shift_data[61] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[61] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[61] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[61] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[61] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[61] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[62] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [62]),
	.C(\macro_inst|controller|serial|shift_data [38]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [62]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~127_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [62]));
defparam \macro_inst|controller|serial|shift_data[62] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[62] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[62] .coord_z = 11;
defparam \macro_inst|controller|serial|shift_data[62] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[62] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[62] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[62] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[62] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[62] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[63] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [39]),
	.C(\macro_inst|controller|sm_pwm|data [63]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [63]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~128_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [63]));
defparam \macro_inst|controller|serial|shift_data[63] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[63] .coord_y = 10;
defparam \macro_inst|controller|serial|shift_data[63] .coord_z = 12;
defparam \macro_inst|controller|serial|shift_data[63] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[63] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[63] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[63] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[63] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[63] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[64] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [40]),
	.C(\macro_inst|controller|sm_pwm|data [64]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [64]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~129_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [64]));
defparam \macro_inst|controller|serial|shift_data[64] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[64] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[64] .coord_z = 12;
defparam \macro_inst|controller|serial|shift_data[64] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[64] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[64] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[64] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[64] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[64] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[65] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [65]),
	.C(\macro_inst|controller|serial|shift_data [41]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [65]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~130_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [65]));
defparam \macro_inst|controller|serial|shift_data[65] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[65] .coord_y = 4;
defparam \macro_inst|controller|serial|shift_data[65] .coord_z = 6;
defparam \macro_inst|controller|serial|shift_data[65] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[65] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[65] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[65] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[65] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[65] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[66] (
	.A(\macro_inst|controller|serial|shift_data [42]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [66]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [66]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~131_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [66]));
defparam \macro_inst|controller|serial|shift_data[66] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[66] .coord_y = 4;
defparam \macro_inst|controller|serial|shift_data[66] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[66] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[66] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[66] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[66] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[66] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[66] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[67] (
	.A(\macro_inst|controller|serial|shift_data [43]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [67]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [67]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~132_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [67]));
defparam \macro_inst|controller|serial|shift_data[67] .coord_x = 17;
defparam \macro_inst|controller|serial|shift_data[67] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[67] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[67] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[67] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[67] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[67] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[67] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[67] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[68] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [68]),
	.C(\macro_inst|controller|serial|shift_data [44]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [68]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~134_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [68]));
defparam \macro_inst|controller|serial|shift_data[68] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[68] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[68] .coord_z = 7;
defparam \macro_inst|controller|serial|shift_data[68] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[68] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[68] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[68] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[68] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[68] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[69] (
	.A(\macro_inst|controller|serial|shift_data [45]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [69]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [69]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~135_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [69]));
defparam \macro_inst|controller|serial|shift_data[69] .coord_x = 14;
defparam \macro_inst|controller|serial|shift_data[69] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[69] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[69] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[69] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[69] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[69] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[69] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[69] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[6] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [6]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [6]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~189_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [6]));
defparam \macro_inst|controller|serial|shift_data[6] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[6] .coord_y = 10;
defparam \macro_inst|controller|serial|shift_data[6] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[6] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[6] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[6] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[70] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [46]),
	.C(\macro_inst|controller|sm_pwm|data [70]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [70]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~136_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [70]));
defparam \macro_inst|controller|serial|shift_data[70] .coord_x = 14;
defparam \macro_inst|controller|serial|shift_data[70] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[70] .coord_z = 4;
defparam \macro_inst|controller|serial|shift_data[70] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[70] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[70] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[70] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[70] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[70] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[71] (
	.A(\macro_inst|controller|serial|shift_data [47]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [71]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [71]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~137_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [71]));
defparam \macro_inst|controller|serial|shift_data[71] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[71] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[71] .coord_z = 14;
defparam \macro_inst|controller|serial|shift_data[71] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[71] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[71] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[71] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[71] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[71] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[72] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [72]),
	.D(\macro_inst|controller|serial|shift_data [48]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [72]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~97_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [72]));
defparam \macro_inst|controller|serial|shift_data[72] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[72] .coord_y = 9;
defparam \macro_inst|controller|serial|shift_data[72] .coord_z = 14;
defparam \macro_inst|controller|serial|shift_data[72] .mask = 16'hAF05;
defparam \macro_inst|controller|serial|shift_data[72] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[72] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[72] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[72] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[72] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[73] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [49]),
	.C(\macro_inst|controller|sm_pwm|data [73]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [73]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~98_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [73]));
defparam \macro_inst|controller|serial|shift_data[73] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[73] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[73] .coord_z = 11;
defparam \macro_inst|controller|serial|shift_data[73] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[73] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[73] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[73] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[73] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[73] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[74] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [50]),
	.C(\macro_inst|controller|sm_pwm|data [74]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [74]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~109_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [74]));
defparam \macro_inst|controller|serial|shift_data[74] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[74] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[74] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[74] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[74] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[74] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[74] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[74] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[74] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[75] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [51]),
	.C(\macro_inst|controller|sm_pwm|data [75]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [75]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~114_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [75]));
defparam \macro_inst|controller|serial|shift_data[75] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[75] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[75] .coord_z = 13;
defparam \macro_inst|controller|serial|shift_data[75] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[75] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[75] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[75] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[75] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[75] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[76] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [76]),
	.C(\macro_inst|controller|serial|shift_data [52]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [76]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~115_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [76]));
defparam \macro_inst|controller|serial|shift_data[76] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[76] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[76] .coord_z = 3;
defparam \macro_inst|controller|serial|shift_data[76] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[76] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[76] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[76] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[76] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[76] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[77] (
	.A(\macro_inst|controller|serial|shift_data [53]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [77]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [77]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~116_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [77]));
defparam \macro_inst|controller|serial|shift_data[77] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[77] .coord_y = 9;
defparam \macro_inst|controller|serial|shift_data[77] .coord_z = 4;
defparam \macro_inst|controller|serial|shift_data[77] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[77] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[77] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[77] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[77] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[77] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[78] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [78]),
	.C(\macro_inst|controller|serial|shift_data [54]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [78]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~117_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [78]));
defparam \macro_inst|controller|serial|shift_data[78] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[78] .coord_y = 10;
defparam \macro_inst|controller|serial|shift_data[78] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[78] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[78] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[78] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[78] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[78] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[78] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[79] (
	.A(\macro_inst|controller|sm_pwm|data [79]),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [55]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [79]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~118_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [79]));
defparam \macro_inst|controller|serial|shift_data[79] .coord_x = 17;
defparam \macro_inst|controller|serial|shift_data[79] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[79] .coord_z = 0;
defparam \macro_inst|controller|serial|shift_data[79] .mask = 16'hF055;
defparam \macro_inst|controller|serial|shift_data[79] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[79] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[79] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[79] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[79] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[7] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [7]),
	.C(vcc),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [7]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~190_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [7]));
defparam \macro_inst|controller|serial|shift_data[7] .coord_x = 17;
defparam \macro_inst|controller|serial|shift_data[7] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[7] .coord_z = 13;
defparam \macro_inst|controller|serial|shift_data[7] .mask = 16'h0033;
defparam \macro_inst|controller|serial|shift_data[7] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[7] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[80] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [80]),
	.D(\macro_inst|controller|serial|shift_data [56]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [80]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~119_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [80]));
defparam \macro_inst|controller|serial|shift_data[80] .coord_x = 11;
defparam \macro_inst|controller|serial|shift_data[80] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[80] .coord_z = 1;
defparam \macro_inst|controller|serial|shift_data[80] .mask = 16'hAF05;
defparam \macro_inst|controller|serial|shift_data[80] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[80] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[80] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[80] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[80] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[81] (
	.A(vcc),
	.B(\macro_inst|controller|serial|state.IDLE~q ),
	.C(\macro_inst|controller|serial|shift_data [57]),
	.D(\macro_inst|controller|sm_pwm|data [81]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [81]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~120_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [81]));
defparam \macro_inst|controller|serial|shift_data[81] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[81] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[81] .coord_z = 1;
defparam \macro_inst|controller|serial|shift_data[81] .mask = 16'hC0F3;
defparam \macro_inst|controller|serial|shift_data[81] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[81] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[81] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[81] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[81] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[82] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [58]),
	.C(\macro_inst|controller|sm_pwm|data [82]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [82]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~99_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [82]));
defparam \macro_inst|controller|serial|shift_data[82] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[82] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[82] .coord_z = 9;
defparam \macro_inst|controller|serial|shift_data[82] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[82] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[82] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[82] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[82] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[82] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[83] (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [59]),
	.D(\macro_inst|controller|sm_pwm|data [83]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [83]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~100_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [83]));
defparam \macro_inst|controller|serial|shift_data[83] .coord_x = 11;
defparam \macro_inst|controller|serial|shift_data[83] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[83] .coord_z = 8;
defparam \macro_inst|controller|serial|shift_data[83] .mask = 16'hA0F5;
defparam \macro_inst|controller|serial|shift_data[83] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[83] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[83] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[83] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[83] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[84] (
	.A(\macro_inst|controller|serial|shift_data [60]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [84]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [84]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~101_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [84]));
defparam \macro_inst|controller|serial|shift_data[84] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[84] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[84] .coord_z = 15;
defparam \macro_inst|controller|serial|shift_data[84] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[84] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[84] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[84] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[84] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[84] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[85] (
	.A(\macro_inst|controller|serial|shift_data [61]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [85]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [85]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~102_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [85]));
defparam \macro_inst|controller|serial|shift_data[85] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[85] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[85] .coord_z = 7;
defparam \macro_inst|controller|serial|shift_data[85] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[85] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[85] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[85] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[85] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[85] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[86] (
	.A(vcc),
	.B(\macro_inst|controller|serial|state.IDLE~q ),
	.C(\macro_inst|controller|serial|shift_data [62]),
	.D(\macro_inst|controller|sm_pwm|data [86]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [86]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X51_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~103_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [86]));
defparam \macro_inst|controller|serial|shift_data[86] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[86] .coord_y = 2;
defparam \macro_inst|controller|serial|shift_data[86] .coord_z = 9;
defparam \macro_inst|controller|serial|shift_data[86] .mask = 16'hC0F3;
defparam \macro_inst|controller|serial|shift_data[86] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[86] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[86] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[86] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[86] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[87] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [63]),
	.C(\macro_inst|controller|sm_pwm|data [87]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [87]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~104_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [87]));
defparam \macro_inst|controller|serial|shift_data[87] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[87] .coord_y = 10;
defparam \macro_inst|controller|serial|shift_data[87] .coord_z = 13;
defparam \macro_inst|controller|serial|shift_data[87] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[87] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[87] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[87] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[87] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[87] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[88] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [64]),
	.C(\macro_inst|controller|sm_pwm|data [88]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [88]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X62_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~105_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [88]));
defparam \macro_inst|controller|serial|shift_data[88] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[88] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[88] .coord_z = 6;
defparam \macro_inst|controller|serial|shift_data[88] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[88] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[88] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[88] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[88] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[88] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[89] (
	.A(\macro_inst|controller|sm_pwm|data [89]),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [65]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [89]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~106_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [89]));
defparam \macro_inst|controller|serial|shift_data[89] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[89] .coord_y = 4;
defparam \macro_inst|controller|serial|shift_data[89] .coord_z = 8;
defparam \macro_inst|controller|serial|shift_data[89] .mask = 16'hF055;
defparam \macro_inst|controller|serial|shift_data[89] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[89] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[89] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[89] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[89] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[8] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|sm_pwm|data [8]),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [8]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~191_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [8]));
defparam \macro_inst|controller|serial|shift_data[8] .coord_x = 11;
defparam \macro_inst|controller|serial|shift_data[8] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[8] .coord_z = 0;
defparam \macro_inst|controller|serial|shift_data[8] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[8] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[8] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[8] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[90] (
	.A(\macro_inst|controller|serial|shift_data [66]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [90]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [90]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~107_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [90]));
defparam \macro_inst|controller|serial|shift_data[90] .coord_x = 15;
defparam \macro_inst|controller|serial|shift_data[90] .coord_y = 4;
defparam \macro_inst|controller|serial|shift_data[90] .coord_z = 10;
defparam \macro_inst|controller|serial|shift_data[90] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[90] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[90] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[90] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[90] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[90] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[91] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [91]),
	.C(\macro_inst|controller|serial|shift_data [67]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [91]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~108_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [91]));
defparam \macro_inst|controller|serial|shift_data[91] .coord_x = 18;
defparam \macro_inst|controller|serial|shift_data[91] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[91] .coord_z = 2;
defparam \macro_inst|controller|serial|shift_data[91] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[91] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[91] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[91] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[91] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[91] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[92] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [68]),
	.C(\macro_inst|controller|sm_pwm|data [92]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [92]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~110_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [92]));
defparam \macro_inst|controller|serial|shift_data[92] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[92] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[92] .coord_z = 6;
defparam \macro_inst|controller|serial|shift_data[92] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[92] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[92] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[92] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[92] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[92] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[93] (
	.A(\macro_inst|controller|sm_pwm|data [93]),
	.B(vcc),
	.C(\macro_inst|controller|serial|shift_data [69]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [93]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~111_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [93]));
defparam \macro_inst|controller|serial|shift_data[93] .coord_x = 14;
defparam \macro_inst|controller|serial|shift_data[93] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[93] .coord_z = 5;
defparam \macro_inst|controller|serial|shift_data[93] .mask = 16'hF055;
defparam \macro_inst|controller|serial|shift_data[93] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[93] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[93] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[93] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[93] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[94] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [94]),
	.C(\macro_inst|controller|serial|shift_data [70]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [94]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~112_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [94]));
defparam \macro_inst|controller|serial|shift_data[94] .coord_x = 14;
defparam \macro_inst|controller|serial|shift_data[94] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[94] .coord_z = 6;
defparam \macro_inst|controller|serial|shift_data[94] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[94] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[94] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[94] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[94] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[94] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[95] (
	.A(\macro_inst|controller|serial|shift_data [71]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [95]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [95]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~113_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [95]));
defparam \macro_inst|controller|serial|shift_data[95] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[95] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[95] .coord_z = 9;
defparam \macro_inst|controller|serial|shift_data[95] .mask = 16'hAA0F;
defparam \macro_inst|controller|serial|shift_data[95] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[95] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[95] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[95] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[95] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[96] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [72]),
	.C(\macro_inst|controller|sm_pwm|data [96]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [96]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X61_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~73_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [96]));
defparam \macro_inst|controller|serial|shift_data[96] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[96] .coord_y = 6;
defparam \macro_inst|controller|serial|shift_data[96] .coord_z = 6;
defparam \macro_inst|controller|serial|shift_data[96] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[96] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[96] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[96] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[96] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[96] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[97] (
	.A(vcc),
	.B(\macro_inst|controller|serial|shift_data [73]),
	.C(\macro_inst|controller|sm_pwm|data [97]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [97]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X52_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X52_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~74_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [97]));
defparam \macro_inst|controller|serial|shift_data[97] .coord_x = 16;
defparam \macro_inst|controller|serial|shift_data[97] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[97] .coord_z = 10;
defparam \macro_inst|controller|serial|shift_data[97] .mask = 16'hCC0F;
defparam \macro_inst|controller|serial|shift_data[97] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[97] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[97] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[97] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[97] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[98] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [98]),
	.C(\macro_inst|controller|serial|shift_data [74]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [98]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X56_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~85_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [98]));
defparam \macro_inst|controller|serial|shift_data[98] .coord_x = 20;
defparam \macro_inst|controller|serial|shift_data[98] .coord_y = 8;
defparam \macro_inst|controller|serial|shift_data[98] .coord_z = 14;
defparam \macro_inst|controller|serial|shift_data[98] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[98] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[98] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[98] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[98] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[98] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[99] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|data [99]),
	.C(\macro_inst|controller|serial|shift_data [75]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [99]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X53_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~90_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [99]));
defparam \macro_inst|controller|serial|shift_data[99] .coord_x = 19;
defparam \macro_inst|controller|serial|shift_data[99] .coord_y = 5;
defparam \macro_inst|controller|serial|shift_data[99] .coord_z = 10;
defparam \macro_inst|controller|serial|shift_data[99] .mask = 16'hF033;
defparam \macro_inst|controller|serial|shift_data[99] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[99] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[99] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[99] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[99] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shift_data[9] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|data [9]),
	.D(\macro_inst|controller|serial|state.IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|shift_data [9]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|shift_data[47]~1_combout_X50_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shift_data~192_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|shift_data [9]));
defparam \macro_inst|controller|serial|shift_data[9] .coord_x = 9;
defparam \macro_inst|controller|serial|shift_data[9] .coord_y = 1;
defparam \macro_inst|controller|serial|shift_data[9] .coord_z = 9;
defparam \macro_inst|controller|serial|shift_data[9] .mask = 16'h000F;
defparam \macro_inst|controller|serial|shift_data[9] .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shift_data[9] .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shift_data[9] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|shi~0 (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|serial|Equal0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|shi~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|shi~0 .coord_x = 7;
defparam \macro_inst|controller|serial|shi~0 .coord_y = 1;
defparam \macro_inst|controller|serial|shi~0 .coord_z = 3;
defparam \macro_inst|controller|serial|shi~0 .mask = 16'h00F0;
defparam \macro_inst|controller|serial|shi~0 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|shi~0 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|shi~0 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|shi~0 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|shi~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|state.IDLE (
	.A(\macro_inst|controller|serial|state.LATCH~q ),
	.B(\macro_inst|controller|serial|state~14_combout ),
	.C(vcc),
	.D(\macro_inst|controller|serial|Equal0~0_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|state.IDLE~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X51_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|state~15_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|state.IDLE~q ));
defparam \macro_inst|controller|serial|state.IDLE .coord_x = 8;
defparam \macro_inst|controller|serial|state.IDLE .coord_y = 1;
defparam \macro_inst|controller|serial|state.IDLE .coord_z = 2;
defparam \macro_inst|controller|serial|state.IDLE .mask = 16'hFC5C;
defparam \macro_inst|controller|serial|state.IDLE .modeMux = 1'b0;
defparam \macro_inst|controller|serial|state.IDLE .FeedbackMux = 1'b1;
defparam \macro_inst|controller|serial|state.IDLE .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|state.IDLE .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|state.IDLE .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|state.LATCH (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|controller|serial|state.SHIFT~q ),
	.D(\macro_inst|controller|serial|Selector4~2_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|state.LATCH~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|Equal0~0_combout_X50_Y1_SIG_INV ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|Selector4~3_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|state.LATCH~q ));
defparam \macro_inst|controller|serial|state.LATCH .coord_x = 7;
defparam \macro_inst|controller|serial|state.LATCH .coord_y = 1;
defparam \macro_inst|controller|serial|state.LATCH .coord_z = 7;
defparam \macro_inst|controller|serial|state.LATCH .mask = 16'hF000;
defparam \macro_inst|controller|serial|state.LATCH .modeMux = 1'b0;
defparam \macro_inst|controller|serial|state.LATCH .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|state.LATCH .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|state.LATCH .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|state.LATCH .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|state.LOAD (
	.A(vcc),
	.B(\macro_inst|controller|serial|Selector2~0_combout ),
	.C(\macro_inst|controller|serial|state~14_combout ),
	.D(\macro_inst|controller|serial|Equal0~0_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|state.LOAD~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X50_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y1_SIG ),
	.SyncReset(SyncReset_X50_Y1_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|controller|serial|state.IDLE~q__SyncLoad_X50_Y1_INV ),
	.LutOut(\macro_inst|controller|serial|state.LOAD~0_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|state.LOAD~q ));
defparam \macro_inst|controller|serial|state.LOAD .coord_x = 7;
defparam \macro_inst|controller|serial|state.LOAD .coord_y = 1;
defparam \macro_inst|controller|serial|state.LOAD .coord_z = 1;
defparam \macro_inst|controller|serial|state.LOAD .mask = 16'hF0CC;
defparam \macro_inst|controller|serial|state.LOAD .modeMux = 1'b0;
defparam \macro_inst|controller|serial|state.LOAD .FeedbackMux = 1'b1;
defparam \macro_inst|controller|serial|state.LOAD .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|state.LOAD .BypassEn = 1'b1;
defparam \macro_inst|controller|serial|state.LOAD .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|state.SHIFT (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|serial|state.LOAD~q ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|state.SHIFT~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|serial|Equal0~0_combout_X50_Y1_SIG_INV ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|state.SHIFT~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|state.SHIFT~q ));
defparam \macro_inst|controller|serial|state.SHIFT .coord_x = 7;
defparam \macro_inst|controller|serial|state.SHIFT .coord_y = 1;
defparam \macro_inst|controller|serial|state.SHIFT .coord_z = 12;
defparam \macro_inst|controller|serial|state.SHIFT .mask = 16'hFF00;
defparam \macro_inst|controller|serial|state.SHIFT .modeMux = 1'b0;
defparam \macro_inst|controller|serial|state.SHIFT .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|state.SHIFT .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|state.SHIFT .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|state.SHIFT .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|state~14 (
	.A(vcc),
	.B(\macro_inst|controller|serialOutputTrigger [1]),
	.C(vcc),
	.D(\macro_inst|controller|serialOutputTrigger [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|state~14_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|state~14 .coord_x = 8;
defparam \macro_inst|controller|serial|state~14 .coord_y = 1;
defparam \macro_inst|controller|serial|state~14 .coord_z = 11;
defparam \macro_inst|controller|serial|state~14 .mask = 16'hFFCC;
defparam \macro_inst|controller|serial|state~14 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|state~14 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|state~14 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|state~14 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|state~14 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sto (
	.A(\macro_inst|controller|serial|state.IDLE~q ),
	.B(\macro_inst|controller|serial|state.LATCH~q ),
	.C(\macro_inst|controller|serial|sto~0_combout ),
	.D(\macro_inst|controller|serial|Equal0~0_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|serial|sto~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X50_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X50_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sto~1_combout ),
	.Cout(),
	.Q(\macro_inst|controller|serial|sto~q ));
defparam \macro_inst|controller|serial|sto .coord_x = 7;
defparam \macro_inst|controller|serial|sto .coord_y = 1;
defparam \macro_inst|controller|serial|sto .coord_z = 4;
defparam \macro_inst|controller|serial|sto .mask = 16'hF0F8;
defparam \macro_inst|controller|serial|sto .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sto .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sto .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sto .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sto .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|serial|sto~0 (
	.A(\macro_inst|controller|serial|sto~q ),
	.B(\macro_inst|controller|serialOutputTrigger [0]),
	.C(\macro_inst|controller|serial|state.IDLE~q ),
	.D(\macro_inst|controller|serialOutputTrigger [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|serial|sto~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|serial|sto~0 .coord_x = 7;
defparam \macro_inst|controller|serial|sto~0 .coord_y = 1;
defparam \macro_inst|controller|serial|sto~0 .coord_z = 14;
defparam \macro_inst|controller|serial|sto~0 .mask = 16'hA0A2;
defparam \macro_inst|controller|serial|sto~0 .modeMux = 1'b0;
defparam \macro_inst|controller|serial|sto~0 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|serial|sto~0 .ShiftMux = 1'b0;
defparam \macro_inst|controller|serial|sto~0 .BypassEn = 1'b0;
defparam \macro_inst|controller|serial|sto~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Add0~14 (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|Add0~13 ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Add0~14_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Add0~14 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Add0~14 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|Add0~14 .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|Add0~14 .mask = 16'h3C3C;
defparam \macro_inst|controller|sm_pwm|Add0~14 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|Add0~14 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Add0~14 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Add0~14 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Add0~14 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~11 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~10_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.C(\macro_inst|ahb_add_reg [4]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~11_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~11 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|Decoder0~11 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~11 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|Decoder0~11 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~11 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~11 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~17 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~15_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~16_combout ),
	.C(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.D(\macro_inst|ahb_add_reg [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~17_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~17 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~17 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|Decoder0~17 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|Decoder0~17 .mask = 16'h0080;
defparam \macro_inst|controller|sm_pwm|Decoder0~17 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~17 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~17 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~17 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~17 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~20 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~18_combout ),
	.C(\macro_inst|ahb_add_reg [6]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~19_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~20_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~20 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~20 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~20 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|Decoder0~20 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~20 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~20 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~20 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~20 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~20 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~21 (
	.A(\macro_inst|ahb_add_reg [6]),
	.B(\macro_inst|ahb_add_reg [5]),
	.C(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.D(\macro_inst|ahb_add_reg [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~21_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~21 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~21 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|Decoder0~21 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|Decoder0~21 .mask = 16'h4000;
defparam \macro_inst|controller|sm_pwm|Decoder0~21 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~21 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~21 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~21 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~21 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~23 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~22_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~12_combout ),
	.C(\macro_inst|ahb_add_reg [6]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~23_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~23 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|Decoder0~23 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|Decoder0~23 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|Decoder0~23 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~23 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~23 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~23 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~23 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~23 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~24 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.B(\macro_inst|ahb_add_reg [6]),
	.C(\macro_inst|controller|sm_pwm|Decoder0~22_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~15_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~24_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~24 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|Decoder0~24 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|Decoder0~24 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|Decoder0~24 .mask = 16'h2000;
defparam \macro_inst|controller|sm_pwm|Decoder0~24 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~24 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~24 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~24 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~24 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~25 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~22_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~18_combout ),
	.C(\macro_inst|ahb_add_reg [6]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~25_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~25 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|Decoder0~25 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|Decoder0~25 .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~25 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~25 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~25 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~25 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~25 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~25 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~26 (
	.A(vcc),
	.B(\macro_inst|ahb_add_reg [5]),
	.C(\macro_inst|ahb_add_reg [6]),
	.D(\macro_inst|controller|sm_pwm|motor_flags[0]~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~26_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~26 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~26 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|Decoder0~26 .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|Decoder0~26 .mask = 16'h3000;
defparam \macro_inst|controller|sm_pwm|Decoder0~26 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~26 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~26 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~26 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~26 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~27 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~8_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~6_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags[0]~3_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~26_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~27_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~27 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~27 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|Decoder0~27 .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|Decoder0~27 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~27 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~27 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~27 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~27 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~27 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~28 (
	.A(\macro_inst|ahb_add_reg [4]),
	.B(\macro_inst|ahb_add_reg [1]),
	.C(\macro_inst|controller|sm_pwm|Decoder0~27_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~28_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~28 .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|Decoder0~28 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|Decoder0~28 .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|Decoder0~28 .mask = 16'h4000;
defparam \macro_inst|controller|sm_pwm|Decoder0~28 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~28 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~28 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~28 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~28 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~29 (
	.A(vcc),
	.B(\macro_inst|ahb_add_reg [5]),
	.C(\macro_inst|ahb_add_reg [1]),
	.D(\macro_inst|ahb_add_reg [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~29_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~29 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|Decoder0~29 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~29 .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|Decoder0~29 .mask = 16'h3000;
defparam \macro_inst|controller|sm_pwm|Decoder0~29 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~29 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~29 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~29 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~29 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~30 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~12_combout ),
	.B(\macro_inst|ahb_add_reg [4]),
	.C(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~29_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~30_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~30 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|Decoder0~30 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|Decoder0~30 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|Decoder0~30 .mask = 16'h2000;
defparam \macro_inst|controller|sm_pwm|Decoder0~30 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~30 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~30 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~30 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~30 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~31 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~27_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~15_combout ),
	.C(\macro_inst|ahb_add_reg [4]),
	.D(\macro_inst|ahb_add_reg [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~31_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~31 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~31 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|Decoder0~31 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|Decoder0~31 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~31 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~31 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~31 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~31 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~31 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~33 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~18_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~32_combout ),
	.C(\macro_inst|ahb_add_reg [1]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~33_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~33 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|Decoder0~33 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|Decoder0~33 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|Decoder0~33 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~33 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~33 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~33 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~33 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~33 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~34 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~13_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~15_combout ),
	.C(\macro_inst|ahb_add_reg [6]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~34_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~34 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~34 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|Decoder0~34 .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|Decoder0~34 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~34 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~34 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~34 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~34 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~34 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~36 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~35_combout ),
	.B(\macro_inst|ahb_add_reg [1]),
	.C(\macro_inst|controller|sm_pwm|Decoder0~4_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~36_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~36 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~36 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|Decoder0~36 .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|Decoder0~36 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~36 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~36 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~36 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~36 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~36 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~37 (
	.A(vcc),
	.B(\macro_inst|ahb_add_reg [1]),
	.C(\macro_inst|ahb_add_reg [5]),
	.D(\macro_inst|ahb_add_reg [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~37_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~37 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~37 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|Decoder0~37 .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~37 .mask = 16'h0C00;
defparam \macro_inst|controller|sm_pwm|Decoder0~37 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~37 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~37 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~37 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~37 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~38 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~12_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~37_combout ),
	.C(\macro_inst|ahb_add_reg [6]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~38_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~38 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~38 .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|Decoder0~38 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|Decoder0~38 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~38 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~38 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~38 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~38 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~38 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~39 (
	.A(\macro_inst|ahb_add_reg [6]),
	.B(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.C(\macro_inst|controller|sm_pwm|Decoder0~15_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~37_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~39_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~39 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|Decoder0~39 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|Decoder0~39 .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|Decoder0~39 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~39 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~39 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~39 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~39 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~39 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~40 (
	.A(\macro_inst|ahb_add_reg [6]),
	.B(\macro_inst|ahb_add_reg [5]),
	.C(\macro_inst|controller|sm_pwm|Decoder0~5_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~40_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~40 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|Decoder0~40 .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|Decoder0~40 .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|Decoder0~40 .mask = 16'h2000;
defparam \macro_inst|controller|sm_pwm|Decoder0~40 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~40 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~40 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~40 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~40 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~42 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~18_combout ),
	.C(\macro_inst|ahb_add_reg [1]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~41_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~42_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~42 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~42 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~42 .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|Decoder0~42 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~42 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~42 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~42 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~42 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~42 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~43 (
	.A(\macro_inst|ahb_add_reg [6]),
	.B(\macro_inst|controller|sm_pwm|Decoder0~37_combout ),
	.C(\macro_inst|controller|sm_pwm|Decoder0~4_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~43_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~43 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~43 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|Decoder0~43 .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~43 .mask = 16'h4000;
defparam \macro_inst|controller|sm_pwm|Decoder0~43 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~43 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~43 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~43 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~43 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~44 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~12_combout ),
	.B(\macro_inst|ahb_add_reg [4]),
	.C(\macro_inst|controller|sm_pwm|Decoder0~10_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~44_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~44 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|Decoder0~44 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~44 .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|Decoder0~44 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~44 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~44 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~44 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~44 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~44 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~45 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~10_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~15_combout ),
	.C(\macro_inst|ahb_add_reg [4]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~45_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~45 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|Decoder0~45 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~45 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|Decoder0~45 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~45 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~45 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~45 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~45 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~45 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~46 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~5_combout ),
	.C(\macro_inst|ahb_add_reg [5]),
	.D(\macro_inst|ahb_add_reg [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~46_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~46 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~46 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|Decoder0~46 .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~46 .mask = 16'h0008;
defparam \macro_inst|controller|sm_pwm|Decoder0~46 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~46 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~46 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~46 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~46 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~47 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~12_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.C(\macro_inst|ahb_add_reg [4]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~16_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~47_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~47 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|Decoder0~47 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~47 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|Decoder0~47 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~47 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~47 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~47 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~47 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~47 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~48 (
	.A(\macro_inst|ahb_add_reg [5]),
	.B(\macro_inst|ahb_add_reg [1]),
	.C(vcc),
	.D(\macro_inst|ahb_add_reg [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~48_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~48 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~48 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|Decoder0~48 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|Decoder0~48 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|Decoder0~48 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~48 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~48 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~48 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~48 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~49 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~48_combout ),
	.B(\macro_inst|ahb_add_reg [6]),
	.C(\macro_inst|controller|sm_pwm|Decoder0~4_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~49_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~49 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~49 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|Decoder0~49 .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|Decoder0~49 .mask = 16'h2000;
defparam \macro_inst|controller|sm_pwm|Decoder0~49 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~49 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~49 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~49 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~49 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~5 (
	.A(\macro_inst|ahb_add_reg [3]),
	.B(\macro_inst|ahb_add_reg [1]),
	.C(\macro_inst|ahb_add_reg [4]),
	.D(\macro_inst|ahb_add_reg [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~5_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~5 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~5 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|Decoder0~5 .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|Decoder0~5 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~5 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~5 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~5 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~5 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~5 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~50 (
	.A(\macro_inst|ahb_add_reg [1]),
	.B(\macro_inst|controller|sm_pwm|Decoder0~12_combout ),
	.C(\macro_inst|controller|sm_pwm|Decoder0~41_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~50_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~50 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~50 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|Decoder0~50 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|Decoder0~50 .mask = 16'h4000;
defparam \macro_inst|controller|sm_pwm|Decoder0~50 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~50 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~50 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~50 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~50 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~52 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~15_combout ),
	.B(\macro_inst|ahb_add_reg [1]),
	.C(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~51_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~52_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~52 .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|Decoder0~52 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|Decoder0~52 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|Decoder0~52 .mask = 16'h2000;
defparam \macro_inst|controller|sm_pwm|Decoder0~52 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~52 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~52 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~52 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~52 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~54 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~53_combout ),
	.B(\macro_inst|ahb_add_reg [4]),
	.C(\macro_inst|controller|sm_pwm|Decoder0~18_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~54_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~54 .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|Decoder0~54 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|Decoder0~54 .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|Decoder0~54 .mask = 16'h2000;
defparam \macro_inst|controller|sm_pwm|Decoder0~54 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~54 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~54 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~54 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~54 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~56 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~55_combout ),
	.C(\macro_inst|ahb_add_reg [1]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~4_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~56_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~56 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~56 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~56 .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~56 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~56 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~56 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~56 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~56 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~56 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~57 (
	.A(\macro_inst|ahb_add_reg [1]),
	.B(\macro_inst|controller|sm_pwm|Decoder0~12_combout ),
	.C(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~55_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~57_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~57 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~57 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~57 .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|Decoder0~57 .mask = 16'h4000;
defparam \macro_inst|controller|sm_pwm|Decoder0~57 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~57 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~57 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~57 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~57 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~58 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~15_combout ),
	.C(\macro_inst|ahb_add_reg [4]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~53_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~58_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~58 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|Decoder0~58 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|Decoder0~58 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|Decoder0~58 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~58 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~58 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~58 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~58 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~58 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~59 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~18_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~53_combout ),
	.C(\macro_inst|ahb_add_reg [4]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~59_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~59 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~59 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|Decoder0~59 .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|Decoder0~59 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~59 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~59 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~59 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~59 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~59 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~6 (
	.A(\macro_inst|controller|sm_pwm|LessThan0~0_combout ),
	.B(\macro_inst|controller|sm_pwm|Equal0~0_combout ),
	.C(\macro_inst|controller|sm_pwm|Equal0~1_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~6_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~6 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~6 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|Decoder0~6 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|Decoder0~6 .mask = 16'h2AAA;
defparam \macro_inst|controller|sm_pwm|Decoder0~6 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~6 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~6 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~6 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~6 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~60 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~48_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.C(\macro_inst|controller|sm_pwm|Decoder0~4_combout ),
	.D(\macro_inst|ahb_add_reg [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~60_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~60 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~60 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|Decoder0~60 .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|Decoder0~60 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~60 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~60 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~60 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~60 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~60 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~61 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~12_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~27_combout ),
	.C(\macro_inst|ahb_add_reg [4]),
	.D(\macro_inst|ahb_add_reg [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~61_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~61 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~61 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|Decoder0~61 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|Decoder0~61 .mask = 16'h0008;
defparam \macro_inst|controller|sm_pwm|Decoder0~61 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~61 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~61 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~61 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~61 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~62 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~32_combout ),
	.C(\macro_inst|ahb_add_reg [1]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~15_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~62_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~62 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|Decoder0~62 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|Decoder0~62 .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~62 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~62 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~62 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~62 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~62 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~62 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~64 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~18_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.C(\macro_inst|ahb_add_reg [4]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~63_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~64_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~64 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~64 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|Decoder0~64 .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|Decoder0~64 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~64 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~64 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~64 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~64 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~64 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~65 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~15_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~41_combout ),
	.C(\macro_inst|ahb_add_reg [1]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~65_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~65 .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|Decoder0~65 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|Decoder0~65 .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~65 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~65 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~65 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~65 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~65 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~65 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~66 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~63_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~4_combout ),
	.C(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.D(\macro_inst|ahb_add_reg [4]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~66_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~66 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~66 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~66 .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|Decoder0~66 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~66 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~66 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~66 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~66 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~66 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~67 (
	.A(\macro_inst|ahb_add_reg [5]),
	.B(\macro_inst|ahb_add_reg [4]),
	.C(vcc),
	.D(\macro_inst|ahb_add_reg [1]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~67_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~67 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~67 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|Decoder0~67 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|Decoder0~67 .mask = 16'h0044;
defparam \macro_inst|controller|sm_pwm|Decoder0~67 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~67 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~67 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~67 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~67 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~68 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~12_combout ),
	.B(\macro_inst|ahb_add_reg [6]),
	.C(\macro_inst|controller|sm_pwm|Decoder0~67_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~68_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~68 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~68 .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|Decoder0~68 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|Decoder0~68 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~68 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~68 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~68 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~68 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~68 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~69 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~15_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~63_combout ),
	.C(\macro_inst|ahb_add_reg [4]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~69_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~69 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|Decoder0~69 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~69 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|Decoder0~69 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~69 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~69 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~69 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~69 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~69 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~70 (
	.A(\macro_inst|ahb_add_reg [4]),
	.B(\macro_inst|ahb_add_reg [1]),
	.C(\macro_inst|controller|sm_pwm|Decoder0~18_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~27_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~70_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~70 .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|Decoder0~70 .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|Decoder0~70 .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~70 .mask = 16'h2000;
defparam \macro_inst|controller|sm_pwm|Decoder0~70 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~70 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~70 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~70 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~70 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~72 (
	.A(\macro_inst|ahb_add_reg [4]),
	.B(\macro_inst|controller|sm_pwm|Decoder0~18_combout ),
	.C(\macro_inst|controller|sm_pwm|Decoder0~71_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~72_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~72 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|Decoder0~72 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|Decoder0~72 .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|Decoder0~72 .mask = 16'h4000;
defparam \macro_inst|controller|sm_pwm|Decoder0~72 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~72 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~72 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~72 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~72 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~73 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~67_combout ),
	.B(\macro_inst|ahb_add_reg [6]),
	.C(\macro_inst|controller|sm_pwm|Decoder0~4_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~73_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~73 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|Decoder0~73 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|Decoder0~73 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|Decoder0~73 .mask = 16'h2000;
defparam \macro_inst|controller|sm_pwm|Decoder0~73 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~73 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~73 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~73 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~73 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~74 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~12_combout ),
	.C(\macro_inst|ahb_add_reg [6]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~67_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~74_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~74 .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|Decoder0~74 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|Decoder0~74 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|Decoder0~74 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~74 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~74 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~74 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~74 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~74 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~76 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~75_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~15_combout ),
	.C(\macro_inst|ahb_add_reg [1]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~76_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~76 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|Decoder0~76 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|Decoder0~76 .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|Decoder0~76 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~76 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~76 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~76 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~76 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~76 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~77 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~75_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~18_combout ),
	.C(\macro_inst|ahb_add_reg [1]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~77_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~77 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|Decoder0~77 .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|Decoder0~77 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|Decoder0~77 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~77 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~77 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~77 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~77 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~77 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~78 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~53_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~4_combout ),
	.C(\macro_inst|ahb_add_reg [4]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~78_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~78 .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~78 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|Decoder0~78 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|Decoder0~78 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~78 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~78 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~78 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~78 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~78 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~79 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~12_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.C(\macro_inst|ahb_add_reg [4]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~53_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~79_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~79 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|Decoder0~79 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|Decoder0~79 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|Decoder0~79 .mask = 16'h0800;
defparam \macro_inst|controller|sm_pwm|Decoder0~79 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~79 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~79 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~79 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~79 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~80 (
	.A(\macro_inst|ahb_add_reg [3]),
	.B(\macro_inst|ahb_add_reg [2]),
	.C(\macro_inst|ahb_add_reg [4]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~21_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~80_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~80 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~80 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|Decoder0~80 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|Decoder0~80 .mask = 16'h1000;
defparam \macro_inst|controller|sm_pwm|Decoder0~80 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~80 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~80 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~80 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~80 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~81 (
	.A(\macro_inst|ahb_add_reg [3]),
	.B(\macro_inst|ahb_add_reg [2]),
	.C(\macro_inst|ahb_add_reg [4]),
	.D(\macro_inst|controller|sm_pwm|Decoder0~21_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~81_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~81 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~81 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|Decoder0~81 .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|Decoder0~81 .mask = 16'h0100;
defparam \macro_inst|controller|sm_pwm|Decoder0~81 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~81 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~81 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~81 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~81 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Decoder0~9 (
	.A(\macro_inst|controller|sm_pwm|motor_flags[0]~3_combout ),
	.B(\macro_inst|controller|sm_pwm|Decoder0~8_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags[0]~5_combout ),
	.D(\macro_inst|controller|sm_pwm|Decoder0~6_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~9_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Decoder0~9 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Decoder0~9 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|Decoder0~9 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|Decoder0~9 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Decoder0~9 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~9 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~9 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~9 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Decoder0~9 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Equal1~0 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Equal1~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Equal1~0 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|Equal1~0 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|Equal1~0 .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|Equal1~0 .mask = 16'h0080;
defparam \macro_inst|controller|sm_pwm|Equal1~0 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Equal1~0 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Equal1~0 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Equal1~0 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Equal1~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|Equal1~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Equal1~1_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|Equal1~1 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|Equal1~1 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|Equal1~1 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|Equal1~1 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|Equal1~1 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Equal1~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Equal1~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|Equal1~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|Equal1~1 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|LessThan10~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[4][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan10~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan10~1 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|LessThan10~1 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|LessThan10~1 .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|LessThan10~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan10~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan10~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan10~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan10~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan10~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan10~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[4][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan10~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan10~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan10~11 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|LessThan10~11 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|LessThan10~11 .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|LessThan10~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan10~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan10~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan10~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan10~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan10~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan12~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[5][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan12~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan12~1 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|LessThan12~1 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan12~1 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|LessThan12~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan12~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan12~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan12~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan12~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan12~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan12~11 (
	.A(\macro_inst|controller|sm_pwm|pwmList[5][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan12~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan12~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan12~11 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|LessThan12~11 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan12~11 .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|LessThan12~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan12~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan12~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan12~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan12~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan12~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan14~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[6][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan14~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan14~1 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan14~1 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan14~1 .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|LessThan14~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan14~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan14~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan14~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan14~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan14~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan14~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[6][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan14~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan14~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan14~11 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan14~11 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan14~11 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|LessThan14~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan14~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan14~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan14~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan14~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan14~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan16~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[7][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan16~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan16~1 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan16~1 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|LessThan16~1 .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|LessThan16~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan16~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan16~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan16~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan16~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan16~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan16~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[7][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan16~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan16~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan16~11 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan16~11 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|LessThan16~11 .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|LessThan16~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan16~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan16~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan16~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan16~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan16~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan18~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[8][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan18~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan18~1 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|LessThan18~1 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|LessThan18~1 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|LessThan18~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan18~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan18~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan18~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan18~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan18~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan18~11 (
	.A(\macro_inst|controller|sm_pwm|pwmList[8][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan18~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan18~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan18~11 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|LessThan18~11 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|LessThan18~11 .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|LessThan18~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan18~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan18~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan18~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan18~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan18~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan20~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[9][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan20~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan20~1 .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|LessThan20~1 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan20~1 .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|LessThan20~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan20~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan20~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan20~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan20~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan20~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan20~11 (
	.A(\macro_inst|controller|sm_pwm|pwmList[9][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan20~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan20~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan20~11 .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|LessThan20~11 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan20~11 .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|LessThan20~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan20~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan20~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan20~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan20~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan20~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan21~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[10][8]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan21~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan21~1 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|LessThan21~1 .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|LessThan21~1 .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|LessThan21~1 .mask = 16'h0044;
defparam \macro_inst|controller|sm_pwm|LessThan21~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan21~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan21~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan21~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan21~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan21~12 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|pwmList[10][14]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan21~11_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan21~12_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan21~12 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|LessThan21~12 .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|LessThan21~12 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|LessThan21~12 .mask = 16'h5F05;
defparam \macro_inst|controller|sm_pwm|LessThan21~12 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan21~12 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan21~12 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan21~12 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan21~12 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|LessThan24~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[11][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan24~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan24~1 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan24~1 .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|LessThan24~1 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|LessThan24~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan24~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan24~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan24~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan24~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan24~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan24~11 (
	.A(\macro_inst|controller|sm_pwm|pwmList[11][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan24~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan24~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan24~11 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan24~11 .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|LessThan24~11 .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|LessThan24~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan24~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan24~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan24~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan24~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan24~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan24~3 (
	.A(\macro_inst|controller|sm_pwm|pwmList[11][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan24~1_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan24~3_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan24~3 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan24~3 .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|LessThan24~3 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|LessThan24~3 .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|LessThan24~3 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan24~3 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan24~3 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan24~3 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan24~3 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan25~3 (
	.A(\macro_inst|controller|sm_pwm|pwmList[12][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan25~1_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan25~3_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan25~3 .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|LessThan25~3 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|LessThan25~3 .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|LessThan25~3 .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|LessThan25~3 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan25~3 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan25~3 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan25~3 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan25~3 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan25~9 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[12][12]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan25~7_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan25~9_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan25~9 .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|LessThan25~9 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|LessThan25~9 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|LessThan25~9 .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|LessThan25~9 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan25~9 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan25~9 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan25~9 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan25~9 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan28~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[13][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan28~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan28~1 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan28~1 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|LessThan28~1 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|LessThan28~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan28~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan28~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan28~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan28~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan28~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan28~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[13][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan28~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan28~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan28~11 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan28~11 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|LessThan28~11 .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|LessThan28~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan28~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan28~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan28~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan28~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan28~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan28~5 (
	.A(\macro_inst|controller|sm_pwm|pwmList[13][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan28~3_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan28~5_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan28~5 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan28~5 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|LessThan28~5 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|LessThan28~5 .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|LessThan28~5 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan28~5 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan28~5 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan28~5 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan28~5 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan2~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[0][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan2~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan2~1 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|LessThan2~1 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|LessThan2~1 .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|LessThan2~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan2~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan2~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan2~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan2~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan2~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan2~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[0][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan2~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan2~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan2~11 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|LessThan2~11 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|LessThan2~11 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|LessThan2~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan2~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan2~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan2~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan2~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan2~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan30~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[14][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan30~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan30~1 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan30~1 .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|LessThan30~1 .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|LessThan30~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan30~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan30~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan30~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan30~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan30~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan30~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[14][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan30~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan30~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan30~11 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan30~11 .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|LessThan30~11 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|LessThan30~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan30~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan30~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan30~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan30~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan30~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan31~12 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|pwmList[15][14]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan31~11_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan31~12_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan31~12 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan31~12 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan31~12 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|LessThan31~12 .mask = 16'h5F05;
defparam \macro_inst|controller|sm_pwm|LessThan31~12 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan31~12 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan31~12 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan31~12 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan31~12 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|LessThan33~12 (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|pwmList[16][14]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan33~11_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan33~12_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan33~12 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan33~12 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|LessThan33~12 .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|LessThan33~12 .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|LessThan33~12 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan33~12 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan33~12 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan33~12 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan33~12 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|LessThan34~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[16][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan34~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan34~1 .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|LessThan34~1 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan34~1 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|LessThan34~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan34~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan34~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan34~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan34~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan34~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan36~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[17][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan36~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan36~1 .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|LessThan36~1 .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|LessThan36~1 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|LessThan36~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan36~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan36~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan36~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan36~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan36~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan36~11 (
	.A(\macro_inst|controller|sm_pwm|pwmList[17][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan36~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan36~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan36~11 .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|LessThan36~11 .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|LessThan36~11 .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|LessThan36~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan36~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan36~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan36~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan36~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan36~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan37~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[18][8]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan37~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan37~1 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan37~1 .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|LessThan37~1 .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|LessThan37~1 .mask = 16'h0044;
defparam \macro_inst|controller|sm_pwm|LessThan37~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan37~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan37~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan37~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan37~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan38~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[18][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan38~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan38~1 .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|LessThan38~1 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|LessThan38~1 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|LessThan38~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan38~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan38~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan38~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan38~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan38~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan38~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[18][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan38~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan38~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan38~11 .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|LessThan38~11 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|LessThan38~11 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|LessThan38~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan38~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan38~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan38~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan38~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan38~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan40~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[19][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan40~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan40~1 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan40~1 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan40~1 .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|LessThan40~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan40~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan40~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan40~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan40~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan40~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan40~11 (
	.A(\macro_inst|controller|sm_pwm|pwmList[19][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan40~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan40~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan40~11 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan40~11 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan40~11 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|LessThan40~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan40~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan40~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan40~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan40~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan40~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan42~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[20][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan42~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan42~1 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan42~1 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|LessThan42~1 .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|LessThan42~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan42~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan42~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan42~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan42~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan42~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan42~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[20][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan42~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan42~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan42~11 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan42~11 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|LessThan42~11 .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|LessThan42~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan42~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan42~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan42~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan42~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan42~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan43~5 (
	.A(\macro_inst|controller|sm_pwm|pwmList[21][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan43~3_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan43~5_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan43~5 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan43~5 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|LessThan43~5 .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|LessThan43~5 .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|LessThan43~5 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan43~5 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan43~5 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan43~5 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan43~5 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan43~9 (
	.A(\macro_inst|controller|sm_pwm|pwmList[21][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan43~7_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan43~9_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan43~9 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan43~9 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|LessThan43~9 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|LessThan43~9 .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|LessThan43~9 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan43~9 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan43~9 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan43~9 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan43~9 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan46~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[22][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan46~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan46~1 .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|LessThan46~1 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|LessThan46~1 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|LessThan46~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan46~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan46~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan46~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan46~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan46~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan46~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[22][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan46~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan46~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan46~11 .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|LessThan46~11 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|LessThan46~11 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|LessThan46~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan46~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan46~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan46~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan46~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan46~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan48~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[23][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan48~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan48~1 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan48~1 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|LessThan48~1 .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|LessThan48~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan48~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan48~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan48~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan48~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan48~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan48~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[23][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan48~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan48~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan48~11 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan48~11 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|LessThan48~11 .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|LessThan48~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan48~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan48~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan48~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan48~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan48~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan50~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[24][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan50~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan50~1 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan50~1 .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|LessThan50~1 .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|LessThan50~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan50~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan50~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan50~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan50~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan50~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan50~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[24][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan50~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan50~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan50~11 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan50~11 .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|LessThan50~11 .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|LessThan50~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan50~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan50~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan50~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan50~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan50~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan52~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[25][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan52~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan52~1 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|LessThan52~1 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|LessThan52~1 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|LessThan52~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan52~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan52~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan52~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan52~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan52~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan52~11 (
	.A(\macro_inst|controller|sm_pwm|pwmList[25][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan52~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan52~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan52~11 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|LessThan52~11 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|LessThan52~11 .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|LessThan52~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan52~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan52~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan52~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan52~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan52~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan54~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[26][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan54~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan54~1 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan54~1 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|LessThan54~1 .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|LessThan54~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan54~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan54~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan54~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan54~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan54~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan54~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[26][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan54~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan54~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan54~11 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan54~11 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|LessThan54~11 .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|LessThan54~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan54~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan54~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan54~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan54~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan54~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan55~11 (
	.A(\macro_inst|controller|sm_pwm|pwmList[27][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan55~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan55~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan55~11 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|LessThan55~11 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan55~11 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|LessThan55~11 .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|LessThan55~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan55~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan55~12 (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[27][14]~q ),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan55~11_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan55~12_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan55~12 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|LessThan55~12 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan55~12 .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|LessThan55~12 .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|LessThan55~12 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan55~12 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~12 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~12 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~12 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|LessThan55~5 (
	.A(\macro_inst|controller|sm_pwm|pwmList[27][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan55~3_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan55~5_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan55~5 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|LessThan55~5 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan55~5 .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|LessThan55~5 .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|LessThan55~5 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan55~5 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~5 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~5 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~5 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan55~7 (
	.A(\macro_inst|controller|sm_pwm|pwmList[27][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan55~5_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan55~7_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan55~7 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|LessThan55~7 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan55~7 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|LessThan55~7 .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|LessThan55~7 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan55~7 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~7 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~7 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~7 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan55~9 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[27][12]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan55~7_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan55~9_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan55~9 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|LessThan55~9 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan55~9 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|LessThan55~9 .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|LessThan55~9 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan55~9 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~9 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~9 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan55~9 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan58~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[28][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan58~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan58~1 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan58~1 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|LessThan58~1 .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|LessThan58~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan58~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan58~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan58~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan58~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan58~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan58~11 (
	.A(\macro_inst|controller|sm_pwm|pwmList[28][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan58~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan58~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan58~11 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan58~11 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|LessThan58~11 .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|LessThan58~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan58~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan58~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan58~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan58~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan58~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan60~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[29][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan60~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan60~1 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan60~1 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|LessThan60~1 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|LessThan60~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan60~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan60~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan60~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan60~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan60~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan60~11 (
	.A(\macro_inst|controller|sm_pwm|pwmList[29][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan60~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan60~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan60~11 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan60~11 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|LessThan60~11 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|LessThan60~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan60~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan60~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan60~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan60~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan60~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan60~12 (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[29][6]~q ),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan60~11_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan60~12_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan60~12 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan60~12 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|LessThan60~12 .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|LessThan60~12 .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|LessThan60~12 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan60~12 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan60~12 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan60~12 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan60~12 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|LessThan60~9 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[29][4]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan60~7_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan60~9_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan60~9 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan60~9 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|LessThan60~9 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|LessThan60~9 .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|LessThan60~9 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan60~9 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan60~9 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan60~9 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan60~9 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan62~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[30][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan62~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan62~1 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan62~1 .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|LessThan62~1 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|LessThan62~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan62~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan62~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan62~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan62~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan62~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan62~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[30][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan62~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan62~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan62~11 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan62~11 .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|LessThan62~11 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|LessThan62~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan62~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan62~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan62~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan62~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan62~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan64~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[31][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan64~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan64~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan64~11 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|LessThan64~11 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|LessThan64~11 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|LessThan64~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan64~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan64~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan64~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan64~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan64~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan66~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[32][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan66~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan66~1 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|LessThan66~1 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|LessThan66~1 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|LessThan66~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan66~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan66~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan66~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan66~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan66~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan66~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[32][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan66~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan66~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan66~11 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|LessThan66~11 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|LessThan66~11 .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|LessThan66~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan66~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan66~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan66~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan66~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan66~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan67~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[33][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan67~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan67~1 .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|LessThan67~1 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|LessThan67~1 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|LessThan67~1 .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|LessThan67~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan67~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan67~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan67~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan67~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan67~9 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[33][12]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan67~7_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan67~9_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan67~9 .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|LessThan67~9 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|LessThan67~9 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|LessThan67~9 .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|LessThan67~9 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan67~9 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan67~9 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan67~9 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan67~9 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan68~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[33][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan68~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan68~1 .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|LessThan68~1 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|LessThan68~1 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|LessThan68~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan68~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan68~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan68~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan68~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan68~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan69~9 (
	.A(\macro_inst|controller|sm_pwm|pwmList[34][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan69~7_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan69~9_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan69~9 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan69~9 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|LessThan69~9 .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|LessThan69~9 .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|LessThan69~9 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan69~9 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan69~9 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan69~9 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan69~9 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan6~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[2][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan6~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan6~1 .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|LessThan6~1 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|LessThan6~1 .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|LessThan6~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan6~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan6~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan6~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan6~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan6~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan70~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[34][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan70~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan70~1 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan70~1 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|LessThan70~1 .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|LessThan70~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan70~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan70~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan70~12 (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[34][6]~q ),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan70~11_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan70~12_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan70~12 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan70~12 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|LessThan70~12 .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|LessThan70~12 .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|LessThan70~12 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan70~12 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~12 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~12 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~12 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|LessThan70~3 (
	.A(\macro_inst|controller|sm_pwm|pwmList[34][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan70~1_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan70~3_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan70~3 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan70~3 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|LessThan70~3 .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|LessThan70~3 .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|LessThan70~3 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan70~3 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~3 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~3 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~3 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan70~5 (
	.A(\macro_inst|controller|sm_pwm|pwmList[34][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan70~3_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan70~5_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan70~5 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan70~5 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|LessThan70~5 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|LessThan70~5 .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|LessThan70~5 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan70~5 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~5 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~5 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~5 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan70~7 (
	.A(\macro_inst|controller|sm_pwm|pwmList[34][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan70~5_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan70~7_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan70~7 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan70~7 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|LessThan70~7 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|LessThan70~7 .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|LessThan70~7 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan70~7 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~7 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~7 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~7 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan70~9 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[34][4]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan70~7_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan70~9_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan70~9 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan70~9 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|LessThan70~9 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|LessThan70~9 .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|LessThan70~9 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan70~9 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~9 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~9 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan70~9 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan72~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[35][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan72~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan72~1 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan72~1 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|LessThan72~1 .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|LessThan72~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan72~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan72~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan72~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan72~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan72~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan72~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[35][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan72~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan72~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan72~11 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|LessThan72~11 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|LessThan72~11 .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|LessThan72~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan72~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan72~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan72~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan72~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan72~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan74~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[36][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan74~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan74~1 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan74~1 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|LessThan74~1 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|LessThan74~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan74~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan74~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan74~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan74~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan74~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan74~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[36][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan74~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan74~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan74~11 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan74~11 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|LessThan74~11 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|LessThan74~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan74~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan74~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan74~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan74~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan74~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan76~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[37][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan76~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan76~1 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan76~1 .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|LessThan76~1 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|LessThan76~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan76~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan76~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan76~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan76~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan76~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan76~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[37][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan76~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan76~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan76~11 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan76~11 .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|LessThan76~11 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|LessThan76~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan76~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan76~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan76~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan76~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan76~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan78~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[38][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan78~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan78~1 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan78~1 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|LessThan78~1 .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|LessThan78~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan78~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan78~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan78~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan78~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan78~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan78~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[38][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan78~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan78~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan78~11 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan78~11 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|LessThan78~11 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|LessThan78~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan78~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan78~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan78~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan78~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan78~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan7~11 (
	.A(\macro_inst|controller|sm_pwm|pwmList[3][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan7~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan7~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan7~11 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan7~11 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|LessThan7~11 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|LessThan7~11 .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|LessThan7~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan7~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan7~12 (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|pwmList[3][14]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan7~11_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan7~12_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan7~12 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan7~12 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|LessThan7~12 .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|LessThan7~12 .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|LessThan7~12 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan7~12 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~12 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~12 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~12 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|LessThan7~3 (
	.A(\macro_inst|controller|sm_pwm|pwmList[3][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan7~1_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan7~3_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan7~3 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan7~3 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|LessThan7~3 .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|LessThan7~3 .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|LessThan7~3 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan7~3 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~3 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~3 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~3 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan7~5 (
	.A(\macro_inst|controller|sm_pwm|pwmList[3][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan7~3_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan7~5_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan7~5 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan7~5 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|LessThan7~5 .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|LessThan7~5 .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|LessThan7~5 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan7~5 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~5 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~5 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~5 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan7~7 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[3][11]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan7~5_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan7~7_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan7~7 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan7~7 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|LessThan7~7 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|LessThan7~7 .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|LessThan7~7 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan7~7 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~7 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~7 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan7~7 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan80~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[39][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan80~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan80~1 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|LessThan80~1 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|LessThan80~1 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|LessThan80~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan80~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan80~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan80~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan80~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan80~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan80~11 (
	.A(\macro_inst|controller|sm_pwm|pwmList[39][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan80~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan80~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan80~11 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|LessThan80~11 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|LessThan80~11 .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|LessThan80~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan80~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan80~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan80~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan80~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan80~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan82~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[40][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan82~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan82~1 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|LessThan82~1 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|LessThan82~1 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|LessThan82~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan82~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan82~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan82~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan82~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan82~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan82~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[40][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan82~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan82~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan82~11 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|LessThan82~11 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|LessThan82~11 .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|LessThan82~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan82~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan82~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan82~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan82~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan82~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan83~12 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|pwmList[41][14]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan83~11_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan83~12_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan83~12 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|LessThan83~12 .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|LessThan83~12 .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|LessThan83~12 .mask = 16'h5F05;
defparam \macro_inst|controller|sm_pwm|LessThan83~12 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan83~12 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan83~12 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan83~12 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan83~12 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|LessThan86~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[42][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan86~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan86~1 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|LessThan86~1 .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|LessThan86~1 .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|LessThan86~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan86~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan86~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan86~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan86~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan86~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan86~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[42][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan86~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan86~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan86~11 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|LessThan86~11 .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|LessThan86~11 .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|LessThan86~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan86~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan86~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan86~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan86~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan86~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan88~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[43][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan88~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan88~1 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|LessThan88~1 .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|LessThan88~1 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|LessThan88~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan88~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan88~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan88~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan88~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan88~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan8~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[3][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan8~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan8~1 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|LessThan8~1 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|LessThan8~1 .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|LessThan8~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan8~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan8~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan8~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan8~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan8~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan8~11 (
	.A(\macro_inst|controller|sm_pwm|pwmList[3][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan8~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan8~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan8~11 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|LessThan8~11 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|LessThan8~11 .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|LessThan8~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan8~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan8~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan8~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan8~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan8~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan90~1 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[44][0]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan90~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan90~1 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan90~1 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|LessThan90~1 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|LessThan90~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan90~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan90~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan90~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan90~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan90~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan90~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[44][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan90~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan90~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan90~11 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan90~11 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|LessThan90~11 .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|LessThan90~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan90~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan90~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan90~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan90~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan90~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan90~7 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[44][3]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan90~5_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan90~7_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan90~7 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|LessThan90~7 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|LessThan90~7 .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|LessThan90~7 .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|LessThan90~7 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan90~7 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan90~7 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan90~7 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan90~7 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan92~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[45][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan92~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan92~1 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan92~1 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|LessThan92~1 .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|LessThan92~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan92~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan92~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan92~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan92~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan92~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan92~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[45][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan92~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan92~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan92~11 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|LessThan92~11 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|LessThan92~11 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|LessThan92~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan92~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan92~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan92~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan92~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan92~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan94~1 (
	.A(\macro_inst|controller|sm_pwm|pwmList[46][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan94~1_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan94~1 .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|LessThan94~1 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|LessThan94~1 .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|LessThan94~1 .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|LessThan94~1 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan94~1 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan94~1 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan94~1 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan94~1 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan94~11 (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[46][5]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan94~9_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan94~11_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan94~11 .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|LessThan94~11 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|LessThan94~11 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|LessThan94~11 .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|LessThan94~11 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan94~11 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan94~11 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan94~11 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan94~11 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan95~5 (
	.A(\macro_inst|controller|sm_pwm|pwmList[47][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan95~3_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan95~5_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan95~5 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|LessThan95~5 .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|LessThan95~5 .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|LessThan95~5 .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|LessThan95~5 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan95~5 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan95~5 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan95~5 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan95~5 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|LessThan95~9 (
	.A(\macro_inst|controller|sm_pwm|pwmList[47][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan95~7_cout ),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan95~9_cout ),
	.Q());
defparam \macro_inst|controller|sm_pwm|LessThan95~9 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|LessThan95~9 .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|LessThan95~9 .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|LessThan95~9 .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|LessThan95~9 .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|LessThan95~9 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan95~9 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan95~9 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|LessThan95~9 .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|data[0] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[0][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan1~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~264_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [0]));
defparam \macro_inst|controller|sm_pwm|data[0] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[0] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[0] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|data[0] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[100] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[9][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan19~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [100]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~138_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [100]));
defparam \macro_inst|controller|sm_pwm|data[100] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data[100] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[100] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[100] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[100] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[100] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[100] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[100] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[100] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[101] (
	.A(\macro_inst|controller|sm_pwm|pwmList[11][15]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|LessThan23~12_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [101]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~139_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [101]));
defparam \macro_inst|controller|sm_pwm|data[101] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[101] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[101] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|data[101] .mask = 16'h2020;
defparam \macro_inst|controller|sm_pwm|data[101] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[101] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[101] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[101] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[101] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[102] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|LessThan27~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[13][15]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [102]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~140_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [102]));
defparam \macro_inst|controller|sm_pwm|data[102] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[102] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[102] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[102] .mask = 16'h3000;
defparam \macro_inst|controller|sm_pwm|data[102] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[102] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[102] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[102] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[102] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[103] (
	.A(\macro_inst|controller|sm_pwm|LessThan31~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[15][15]~q ),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [103]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y5_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~141_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [103]));
defparam \macro_inst|controller|sm_pwm|data[103] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[103] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|data[103] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[103] .mask = 16'h0088;
defparam \macro_inst|controller|sm_pwm|data[103] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[103] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[103] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[103] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[103] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[104] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[17][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan35~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [104]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~142_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [104]));
defparam \macro_inst|controller|sm_pwm|data[104] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|data[104] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data[104] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|data[104] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[104] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[104] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[104] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[104] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[104] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[105] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|pwmList[19][15]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan39~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [105]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~143_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [105]));
defparam \macro_inst|controller|sm_pwm|data[105] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[105] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[105] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|data[105] .mask = 16'h3000;
defparam \macro_inst|controller|sm_pwm|data[105] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[105] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[105] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[105] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[105] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[106] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|LessThan43~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[21][15]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [106]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~122_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [106]));
defparam \macro_inst|controller|sm_pwm|data[106] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[106] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|data[106] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|data[106] .mask = 16'h5000;
defparam \macro_inst|controller|sm_pwm|data[106] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[106] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[106] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[106] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[106] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[107] (
	.A(\macro_inst|controller|sm_pwm|pwmList[23][15]~q ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|LessThan47~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [107]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~123_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [107]));
defparam \macro_inst|controller|sm_pwm|data[107] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[107] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[107] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[107] .mask = 16'h00A0;
defparam \macro_inst|controller|sm_pwm|data[107] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[107] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[107] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[107] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[107] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[108] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|pwmList[25][15]~q ),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|LessThan51~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [108]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~124_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [108]));
defparam \macro_inst|controller|sm_pwm|data[108] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[108] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data[108] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[108] .mask = 16'h4400;
defparam \macro_inst|controller|sm_pwm|data[108] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[108] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[108] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[108] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[108] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[109] (
	.A(\macro_inst|controller|sm_pwm|LessThan55~12_combout ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmList[27][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [109]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~125_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [109]));
defparam \macro_inst|controller|sm_pwm|data[109] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[109] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data[109] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[109] .mask = 16'h00A0;
defparam \macro_inst|controller|sm_pwm|data[109] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[109] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[109] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[109] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[109] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[10] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|pwmList[20][15]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan41~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [10]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X54_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~266_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [10]));
defparam \macro_inst|controller|sm_pwm|data[10] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[10] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data[10] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[10] .mask = 16'h3000;
defparam \macro_inst|controller|sm_pwm|data[10] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[10] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[10] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[110] (
	.A(\macro_inst|controller|sm_pwm|LessThan59~12_combout ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmList[29][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [110]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~126_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [110]));
defparam \macro_inst|controller|sm_pwm|data[110] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[110] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[110] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|data[110] .mask = 16'h00A0;
defparam \macro_inst|controller|sm_pwm|data[110] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[110] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[110] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[110] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[110] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[111] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[31][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan63~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [111]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~127_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [111]));
defparam \macro_inst|controller|sm_pwm|data[111] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[111] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|data[111] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[111] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[111] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[111] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[111] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[111] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[111] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[112] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|LessThan67~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[33][15]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [112]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~128_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [112]));
defparam \macro_inst|controller|sm_pwm|data[112] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data[112] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data[112] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data[112] .mask = 16'h5000;
defparam \macro_inst|controller|sm_pwm|data[112] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[112] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[112] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[112] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[112] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[113] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|pwmList[35][15]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan71~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [113]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~129_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [113]));
defparam \macro_inst|controller|sm_pwm|data[113] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[113] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data[113] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[113] .mask = 16'h3000;
defparam \macro_inst|controller|sm_pwm|data[113] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[113] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[113] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[113] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[113] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[114] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan75~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[37][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [114]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y5_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~130_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [114]));
defparam \macro_inst|controller|sm_pwm|data[114] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[114] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data[114] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|data[114] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[114] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[114] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[114] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[114] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[114] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[115] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan79~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[39][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [115]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y8_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~131_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [115]));
defparam \macro_inst|controller|sm_pwm|data[115] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[115] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[115] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[115] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[115] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[115] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[115] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[115] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[115] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[116] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|pwmList[41][15]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan83~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [116]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~133_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [116]));
defparam \macro_inst|controller|sm_pwm|data[116] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[116] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|data[116] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[116] .mask = 16'h3000;
defparam \macro_inst|controller|sm_pwm|data[116] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[116] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[116] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[116] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[116] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[117] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan87~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[43][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [117]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~134_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [117]));
defparam \macro_inst|controller|sm_pwm|data[117] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[117] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[117] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[117] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[117] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[117] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[117] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[117] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[117] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[118] (
	.A(\macro_inst|controller|sm_pwm|LessThan91~12_combout ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|pwmList[45][15]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [118]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~135_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [118]));
defparam \macro_inst|controller|sm_pwm|data[118] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[118] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[118] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|data[118] .mask = 16'h0A00;
defparam \macro_inst|controller|sm_pwm|data[118] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[118] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[118] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[118] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[118] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[119] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[47][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan95~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [119]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X60_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~136_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [119]));
defparam \macro_inst|controller|sm_pwm|data[119] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[119] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data[119] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|data[119] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[119] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[119] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[119] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[119] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[119] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[11] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|LessThan45~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[22][15]~q ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [11]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~267_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [11]));
defparam \macro_inst|controller|sm_pwm|data[11] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|data[11] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[11] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|data[11] .mask = 16'h4040;
defparam \macro_inst|controller|sm_pwm|data[11] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[11] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[11] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[120] (
	.A(\macro_inst|controller|sm_pwm|LessThan3~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~72_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [120]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~73_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [120]));
defparam \macro_inst|controller|sm_pwm|data[120] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[120] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[120] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|data[120] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[120] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[120] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[120] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[120] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[120] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[121] (
	.A(\macro_inst|controller|sm_pwm|LessThan7~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|data~74_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [121]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X60_Y6_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~75_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [121]));
defparam \macro_inst|controller|sm_pwm|data[121] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[121] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|data[121] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|data[121] .mask = 16'h000E;
defparam \macro_inst|controller|sm_pwm|data[121] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[121] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[121] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[121] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[121] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[122] (
	.A(\macro_inst|controller|sm_pwm|data~96_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan11~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [122]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~97_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [122]));
defparam \macro_inst|controller|sm_pwm|data[122] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[122] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[122] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[122] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[122] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[122] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[122] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[122] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[122] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[123] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|data~106_combout ),
	.C(\macro_inst|controller|sm_pwm|LessThan15~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [123]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X60_Y6_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~107_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [123]));
defparam \macro_inst|controller|sm_pwm|data[123] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[123] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|data[123] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|data[123] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[123] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[123] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[123] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[123] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[123] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[124] (
	.A(\macro_inst|controller|sm_pwm|data~108_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|LessThan19~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [124]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~109_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [124]));
defparam \macro_inst|controller|sm_pwm|data[124] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data[124] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[124] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[124] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[124] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[124] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[124] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[124] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[124] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[125] (
	.A(\macro_inst|controller|sm_pwm|LessThan23~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~110_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [125]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~111_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [125]));
defparam \macro_inst|controller|sm_pwm|data[125] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[125] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[125] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|data[125] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[125] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[125] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[125] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[125] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[125] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[126] (
	.A(\macro_inst|controller|sm_pwm|data~112_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|LessThan27~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [126]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~113_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [126]));
defparam \macro_inst|controller|sm_pwm|data[126] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[126] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[126] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|data[126] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[126] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[126] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[126] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[126] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[126] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[127] (
	.A(\macro_inst|controller|sm_pwm|data~114_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|LessThan31~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [127]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y8_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~115_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [127]));
defparam \macro_inst|controller|sm_pwm|data[127] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[127] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[127] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|data[127] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[127] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[127] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[127] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[127] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[127] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[128] (
	.A(\macro_inst|controller|sm_pwm|data~116_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan36~12_combout ),
	.C(\macro_inst|controller|sm_pwm|LessThan35~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [128]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~117_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [128]));
defparam \macro_inst|controller|sm_pwm|data[128] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|data[128] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data[128] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[128] .mask = 16'h4450;
defparam \macro_inst|controller|sm_pwm|data[128] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[128] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[128] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[128] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[128] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[129] (
	.A(\macro_inst|controller|sm_pwm|LessThan39~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|data~118_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [129]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~119_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [129]));
defparam \macro_inst|controller|sm_pwm|data[129] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[129] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[129] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[129] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[129] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[129] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[129] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[129] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[129] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[12] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[24][15]~q ),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|LessThan49~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [12]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~268_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [12]));
defparam \macro_inst|controller|sm_pwm|data[12] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[12] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|data[12] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|data[12] .mask = 16'h0C00;
defparam \macro_inst|controller|sm_pwm|data[12] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[12] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[12] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[130] (
	.A(\macro_inst|controller|sm_pwm|LessThan43~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~76_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [130]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~77_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [130]));
defparam \macro_inst|controller|sm_pwm|data[130] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[130] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|data[130] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[130] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[130] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[130] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[130] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[130] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[130] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[131] (
	.A(\macro_inst|controller|sm_pwm|LessThan47~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|data~78_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [131]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~79_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [131]));
defparam \macro_inst|controller|sm_pwm|data[131] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[131] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[131] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[131] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[131] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[131] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[131] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[131] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[131] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[132] (
	.A(\macro_inst|controller|sm_pwm|data~80_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|LessThan51~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [132]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~81_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [132]));
defparam \macro_inst|controller|sm_pwm|data[132] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[132] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data[132] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[132] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[132] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[132] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[132] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[132] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[132] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[133] (
	.A(\macro_inst|controller|sm_pwm|LessThan55~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~82_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [133]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y8_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~83_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [133]));
defparam \macro_inst|controller|sm_pwm|data[133] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[133] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[133] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[133] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[133] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[133] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[133] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[133] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[133] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[134] (
	.A(\macro_inst|controller|sm_pwm|data~84_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan59~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [134]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~85_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [134]));
defparam \macro_inst|controller|sm_pwm|data[134] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[134] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[134] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[134] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[134] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[134] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[134] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[134] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[134] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[135] (
	.A(\macro_inst|controller|sm_pwm|LessThan63~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~86_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [135]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~87_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [135]));
defparam \macro_inst|controller|sm_pwm|data[135] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[135] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|data[135] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|data[135] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[135] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[135] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[135] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[135] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[135] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[136] (
	.A(\macro_inst|controller|sm_pwm|data~88_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|LessThan67~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [136]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~89_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [136]));
defparam \macro_inst|controller|sm_pwm|data[136] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data[136] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data[136] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[136] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[136] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[136] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[136] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[136] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[136] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[137] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|LessThan71~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|data~90_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [137]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~91_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [137]));
defparam \macro_inst|controller|sm_pwm|data[137] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[137] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data[137] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|data[137] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[137] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[137] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[137] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[137] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[137] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[138] (
	.A(\macro_inst|controller|sm_pwm|data~92_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan75~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [138]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y5_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~93_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [138]));
defparam \macro_inst|controller|sm_pwm|data[138] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[138] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data[138] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data[138] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[138] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[138] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[138] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[138] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[138] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[139] (
	.A(\macro_inst|controller|sm_pwm|LessThan79~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|data~94_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [139]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y8_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~95_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [139]));
defparam \macro_inst|controller|sm_pwm|data[139] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[139] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[139] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[139] .mask = 16'h0302;
defparam \macro_inst|controller|sm_pwm|data[139] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[139] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[139] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[139] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[139] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[13] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[26][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan53~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [13]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y6_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~269_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [13]));
defparam \macro_inst|controller|sm_pwm|data[13] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[13] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[13] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[13] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[13] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[13] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[13] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[140] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|data~98_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|LessThan83~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [140]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~99_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [140]));
defparam \macro_inst|controller|sm_pwm|data[140] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[140] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|data[140] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|data[140] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[140] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[140] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[140] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[140] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[140] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[141] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|data~100_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|LessThan87~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [141]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~101_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [141]));
defparam \macro_inst|controller|sm_pwm|data[141] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data[141] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[141] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|data[141] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[141] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[141] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[141] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[141] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[141] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[142] (
	.A(\macro_inst|controller|sm_pwm|LessThan91~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|data~102_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [142]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~103_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [142]));
defparam \macro_inst|controller|sm_pwm|data[142] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[142] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[142] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data[142] .mask = 16'h0302;
defparam \macro_inst|controller|sm_pwm|data[142] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[142] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[142] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[142] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[142] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[143] (
	.A(\macro_inst|controller|sm_pwm|data~104_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan95~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [143]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X60_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~105_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [143]));
defparam \macro_inst|controller|sm_pwm|data[143] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[143] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data[143] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|data[143] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[143] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[143] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[143] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[143] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[143] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[144] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|data~24_combout ),
	.D(\macro_inst|controller|sm_pwm|LessThan4~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [144]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~25_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [144]));
defparam \macro_inst|controller|sm_pwm|data[144] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[144] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[144] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|data[144] .mask = 16'h0302;
defparam \macro_inst|controller|sm_pwm|data[144] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[144] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[144] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[144] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[144] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[145] (
	.A(\macro_inst|controller|sm_pwm|data~26_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|LessThan8~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [145]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~27_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [145]));
defparam \macro_inst|controller|sm_pwm|data[145] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[145] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[145] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[145] .mask = 16'h0504;
defparam \macro_inst|controller|sm_pwm|data[145] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[145] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[145] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[145] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[145] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[146] (
	.A(\macro_inst|controller|sm_pwm|LessThan12~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~48_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [146]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y10_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~49_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [146]));
defparam \macro_inst|controller|sm_pwm|data[146] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[146] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[146] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[146] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[146] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[146] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[146] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[146] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[146] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[147] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|LessThan16~12_combout ),
	.C(\macro_inst|controller|sm_pwm|data~58_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [147]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y10_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~59_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [147]));
defparam \macro_inst|controller|sm_pwm|data[147] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[147] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[147] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[147] .mask = 16'h000E;
defparam \macro_inst|controller|sm_pwm|data[147] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[147] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[147] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[147] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[147] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[148] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|LessThan20~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|data~60_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [148]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~61_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [148]));
defparam \macro_inst|controller|sm_pwm|data[148] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data[148] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[148] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[148] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[148] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[148] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[148] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[148] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[148] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[149] (
	.A(\macro_inst|controller|sm_pwm|data~62_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|LessThan24~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [149]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~63_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [149]));
defparam \macro_inst|controller|sm_pwm|data[149] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[149] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[149] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|data[149] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[149] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[149] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[149] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[149] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[149] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[14] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|LessThan57~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[28][15]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [14]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~270_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [14]));
defparam \macro_inst|controller|sm_pwm|data[14] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[14] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[14] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|data[14] .mask = 16'h5000;
defparam \macro_inst|controller|sm_pwm|data[14] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[14] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[150] (
	.A(\macro_inst|controller|sm_pwm|LessThan27~12_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan28~12_combout ),
	.C(\macro_inst|controller|sm_pwm|data~64_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [150]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~65_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [150]));
defparam \macro_inst|controller|sm_pwm|data[150] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[150] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[150] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|data[150] .mask = 16'h0A0C;
defparam \macro_inst|controller|sm_pwm|data[150] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[150] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[150] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[150] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[150] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[151] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|LessThan32~12_combout ),
	.C(\macro_inst|controller|sm_pwm|data~66_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [151]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~67_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [151]));
defparam \macro_inst|controller|sm_pwm|data[151] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[151] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[151] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|data[151] .mask = 16'h0504;
defparam \macro_inst|controller|sm_pwm|data[151] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[151] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[151] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[151] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[151] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[152] (
	.A(\macro_inst|controller|sm_pwm|data~68_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan36~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [152]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~69_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [152]));
defparam \macro_inst|controller|sm_pwm|data[152] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|data[152] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data[152] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[152] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[152] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[152] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[152] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[152] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[152] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[153] (
	.A(\macro_inst|controller|sm_pwm|LessThan40~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~70_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [153]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~71_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [153]));
defparam \macro_inst|controller|sm_pwm|data[153] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[153] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[153] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[153] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[153] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[153] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[153] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[153] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[153] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[154] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|data~28_combout ),
	.C(\macro_inst|controller|sm_pwm|LessThan44~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [154]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~29_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [154]));
defparam \macro_inst|controller|sm_pwm|data[154] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[154] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|data[154] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|data[154] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[154] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[154] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[154] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[154] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[154] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[155] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|LessThan48~12_combout ),
	.C(\macro_inst|controller|sm_pwm|data~30_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [155]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~31_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [155]));
defparam \macro_inst|controller|sm_pwm|data[155] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[155] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[155] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data[155] .mask = 16'h000E;
defparam \macro_inst|controller|sm_pwm|data[155] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[155] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[155] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[155] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[155] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[156] (
	.A(\macro_inst|controller|sm_pwm|LessThan51~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|data~32_combout ),
	.D(\macro_inst|controller|sm_pwm|LessThan52~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [156]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~33_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [156]));
defparam \macro_inst|controller|sm_pwm|data[156] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[156] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data[156] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[156] .mask = 16'h0B08;
defparam \macro_inst|controller|sm_pwm|data[156] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[156] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[156] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[156] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[156] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[157] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|LessThan56~12_combout ),
	.D(\macro_inst|controller|sm_pwm|data~34_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [157]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~35_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [157]));
defparam \macro_inst|controller|sm_pwm|data[157] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[157] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[157] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|data[157] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[157] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[157] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[157] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[157] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[157] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[158] (
	.A(\macro_inst|controller|sm_pwm|data~36_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|LessThan60~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [158]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~37_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [158]));
defparam \macro_inst|controller|sm_pwm|data[158] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[158] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[158] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[158] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[158] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[158] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[158] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[158] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[158] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[159] (
	.A(\macro_inst|controller|sm_pwm|data~38_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan64~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [159]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~39_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [159]));
defparam \macro_inst|controller|sm_pwm|data[159] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[159] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|data[159] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|data[159] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[159] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[159] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[159] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[159] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[159] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[30][15]~q ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|LessThan61~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [15]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~271_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [15]));
defparam \macro_inst|controller|sm_pwm|data[15] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[15] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|data[15] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|data[15] .mask = 16'h00A0;
defparam \macro_inst|controller|sm_pwm|data[15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[15] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[160] (
	.A(\macro_inst|controller|sm_pwm|data~40_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan68~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [160]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~41_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [160]));
defparam \macro_inst|controller|sm_pwm|data[160] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data[160] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data[160] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|data[160] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[160] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[160] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[160] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[160] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[160] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[161] (
	.A(\macro_inst|controller|sm_pwm|data~42_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan72~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [161]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~43_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [161]));
defparam \macro_inst|controller|sm_pwm|data[161] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[161] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data[161] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|data[161] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[161] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[161] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[161] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[161] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[161] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[162] (
	.A(\macro_inst|controller|sm_pwm|data~44_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan76~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [162]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y5_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~45_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [162]));
defparam \macro_inst|controller|sm_pwm|data[162] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[162] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data[162] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|data[162] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[162] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[162] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[162] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[162] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[162] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[163] (
	.A(\macro_inst|controller|sm_pwm|data~46_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|LessThan80~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [163]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y8_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~47_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [163]));
defparam \macro_inst|controller|sm_pwm|data[163] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[163] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[163] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|data[163] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[163] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[163] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[163] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[163] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[163] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[164] (
	.A(\macro_inst|controller|sm_pwm|LessThan84~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|data~50_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [164]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~51_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [164]));
defparam \macro_inst|controller|sm_pwm|data[164] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[164] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|data[164] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[164] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[164] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[164] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[164] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[164] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[164] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[165] (
	.A(\macro_inst|controller|sm_pwm|LessThan88~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~52_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [165]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~53_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [165]));
defparam \macro_inst|controller|sm_pwm|data[165] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[165] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[165] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|data[165] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[165] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[165] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[165] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[165] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[165] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[166] (
	.A(\macro_inst|controller|sm_pwm|data~54_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|LessThan92~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [166]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~55_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [166]));
defparam \macro_inst|controller|sm_pwm|data[166] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[166] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[166] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|data[166] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[166] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[166] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[166] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[166] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[166] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[167] (
	.A(\macro_inst|controller|sm_pwm|data~56_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan96~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [167]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X60_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~57_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [167]));
defparam \macro_inst|controller|sm_pwm|data[167] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[167] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data[167] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data[167] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[167] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[167] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[167] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[167] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[167] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[168] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|pwmList[1][7]~q ),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|LessThan4~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [168]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~0_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [168]));
defparam \macro_inst|controller|sm_pwm|data[168] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[168] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data[168] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|data[168] .mask = 16'h1100;
defparam \macro_inst|controller|sm_pwm|data[168] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[168] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[168] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[168] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[168] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[169] (
	.A(\macro_inst|controller|sm_pwm|pwmList[3][7]~q ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|LessThan8~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [169]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X60_Y6_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~1_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [169]));
defparam \macro_inst|controller|sm_pwm|data[169] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[169] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|data[169] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[169] .mask = 16'h0500;
defparam \macro_inst|controller|sm_pwm|data[169] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[169] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[169] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[169] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[169] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[16] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[32][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan65~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [16]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~272_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [16]));
defparam \macro_inst|controller|sm_pwm|data[16] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[16] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|data[16] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[16] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[16] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[16] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[16] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[16] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[16] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[170] (
	.A(\macro_inst|controller|sm_pwm|LessThan12~12_combout ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|pwmList[5][7]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [170]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y10_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [170]));
defparam \macro_inst|controller|sm_pwm|data[170] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[170] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[170] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[170] .mask = 16'h000A;
defparam \macro_inst|controller|sm_pwm|data[170] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[170] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[170] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[170] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[170] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[171] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmList[7][7]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan16~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [171]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y10_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~17_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [171]));
defparam \macro_inst|controller|sm_pwm|data[171] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[171] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[171] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data[171] .mask = 16'h0500;
defparam \macro_inst|controller|sm_pwm|data[171] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[171] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[171] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[171] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[171] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[172] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan20~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[9][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [172]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~18_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [172]));
defparam \macro_inst|controller|sm_pwm|data[172] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data[172] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[172] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|data[172] .mask = 16'h000C;
defparam \macro_inst|controller|sm_pwm|data[172] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[172] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[172] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[172] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[172] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[173] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[11][7]~q ),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|LessThan24~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [173]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~19_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [173]));
defparam \macro_inst|controller|sm_pwm|data[173] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[173] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[173] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|data[173] .mask = 16'h0300;
defparam \macro_inst|controller|sm_pwm|data[173] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[173] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[173] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[173] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[173] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[174] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|pwmList[13][7]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan28~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [174]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~20_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [174]));
defparam \macro_inst|controller|sm_pwm|data[174] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[174] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[174] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[174] .mask = 16'h0300;
defparam \macro_inst|controller|sm_pwm|data[174] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[174] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[174] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[174] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[174] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[175] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|pwmList[15][7]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan32~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [175]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~21_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [175]));
defparam \macro_inst|controller|sm_pwm|data[175] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[175] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[175] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[175] .mask = 16'h0300;
defparam \macro_inst|controller|sm_pwm|data[175] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[175] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[175] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[175] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[175] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[176] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan36~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|pwmList[17][7]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [176]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~22_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [176]));
defparam \macro_inst|controller|sm_pwm|data[176] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|data[176] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data[176] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[176] .mask = 16'h000C;
defparam \macro_inst|controller|sm_pwm|data[176] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[176] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[176] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[176] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[176] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[177] (
	.A(\macro_inst|controller|sm_pwm|pwmList[19][7]~q ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|LessThan40~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [177]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~23_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [177]));
defparam \macro_inst|controller|sm_pwm|data[177] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[177] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[177] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|data[177] .mask = 16'h0050;
defparam \macro_inst|controller|sm_pwm|data[177] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[177] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[177] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[177] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[177] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[178] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmList[21][7]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan44~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [178]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~2_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [178]));
defparam \macro_inst|controller|sm_pwm|data[178] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[178] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|data[178] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[178] .mask = 16'h0500;
defparam \macro_inst|controller|sm_pwm|data[178] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[178] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[178] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[178] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[178] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[179] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|LessThan48~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[23][7]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [179]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~3_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [179]));
defparam \macro_inst|controller|sm_pwm|data[179] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[179] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[179] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|data[179] .mask = 16'h0030;
defparam \macro_inst|controller|sm_pwm|data[179] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[179] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[179] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[179] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[179] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[17] (
	.A(\macro_inst|controller|sm_pwm|LessThan69~12_combout ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmList[34][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [17]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~273_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [17]));
defparam \macro_inst|controller|sm_pwm|data[17] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[17] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data[17] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|data[17] .mask = 16'h00A0;
defparam \macro_inst|controller|sm_pwm|data[17] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[17] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[17] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[17] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[17] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[180] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmList[25][7]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan52~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [180]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~4_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [180]));
defparam \macro_inst|controller|sm_pwm|data[180] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[180] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data[180] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[180] .mask = 16'h0500;
defparam \macro_inst|controller|sm_pwm|data[180] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[180] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[180] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[180] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[180] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[181] (
	.A(\macro_inst|controller|sm_pwm|LessThan56~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|pwmList[27][7]~q ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [181]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~5_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [181]));
defparam \macro_inst|controller|sm_pwm|data[181] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[181] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|data[181] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|data[181] .mask = 16'h0202;
defparam \macro_inst|controller|sm_pwm|data[181] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[181] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[181] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[181] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[181] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[182] (
	.A(\macro_inst|controller|sm_pwm|pwmList[29][7]~q ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|LessThan60~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [182]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~6_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [182]));
defparam \macro_inst|controller|sm_pwm|data[182] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[182] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data[182] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|data[182] .mask = 16'h0050;
defparam \macro_inst|controller|sm_pwm|data[182] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[182] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[182] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[182] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[182] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[183] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan64~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[31][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [183]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~7_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [183]));
defparam \macro_inst|controller|sm_pwm|data[183] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[183] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|data[183] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|data[183] .mask = 16'h000C;
defparam \macro_inst|controller|sm_pwm|data[183] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[183] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[183] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[183] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[183] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[184] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan68~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[33][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [184]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~8_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [184]));
defparam \macro_inst|controller|sm_pwm|data[184] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data[184] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data[184] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|data[184] .mask = 16'h000C;
defparam \macro_inst|controller|sm_pwm|data[184] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[184] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[184] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[184] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[184] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[185] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan72~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[35][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [185]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~9_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [185]));
defparam \macro_inst|controller|sm_pwm|data[185] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[185] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data[185] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|data[185] .mask = 16'h000C;
defparam \macro_inst|controller|sm_pwm|data[185] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[185] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[185] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[185] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[185] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[186] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[37][7]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan76~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [186]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y5_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~10_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [186]));
defparam \macro_inst|controller|sm_pwm|data[186] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[186] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data[186] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|data[186] .mask = 16'h0030;
defparam \macro_inst|controller|sm_pwm|data[186] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[186] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[186] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[186] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[186] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[187] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|LessThan80~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[39][7]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [187]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y8_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~11_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [187]));
defparam \macro_inst|controller|sm_pwm|data[187] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[187] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[187] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|data[187] .mask = 16'h0030;
defparam \macro_inst|controller|sm_pwm|data[187] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[187] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[187] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[187] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[187] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[188] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmList[41][7]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan84~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [188]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X60_Y6_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~13_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [188]));
defparam \macro_inst|controller|sm_pwm|data[188] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[188] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|data[188] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|data[188] .mask = 16'h0500;
defparam \macro_inst|controller|sm_pwm|data[188] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[188] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[188] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[188] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[188] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[189] (
	.A(\macro_inst|controller|sm_pwm|pwmList[43][7]~q ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|LessThan88~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [189]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y10_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~14_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [189]));
defparam \macro_inst|controller|sm_pwm|data[189] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[189] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[189] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[189] .mask = 16'h0500;
defparam \macro_inst|controller|sm_pwm|data[189] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[189] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[189] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[189] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[189] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[18] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|pwmList[36][15]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan73~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [18]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~274_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [18]));
defparam \macro_inst|controller|sm_pwm|data[18] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[18] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[18] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[18] .mask = 16'h3000;
defparam \macro_inst|controller|sm_pwm|data[18] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[18] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[18] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[18] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[18] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[190] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|pwmList[45][7]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan92~12_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [190]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~15_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [190]));
defparam \macro_inst|controller|sm_pwm|data[190] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[190] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[190] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[190] .mask = 16'h1010;
defparam \macro_inst|controller|sm_pwm|data[190] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[190] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[190] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[190] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[190] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[191] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan96~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[47][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [191]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X60_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~16_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [191]));
defparam \macro_inst|controller|sm_pwm|data[191] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[191] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data[191] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[191] .mask = 16'h000C;
defparam \macro_inst|controller|sm_pwm|data[191] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[191] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[191] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[191] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[191] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[19] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[38][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan77~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [19]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y5_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~275_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [19]));
defparam \macro_inst|controller|sm_pwm|data[19] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[19] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|data[19] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[19] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[19] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[19] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[19] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[19] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[19] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[1] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[2][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan5~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y10_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~265_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [1]));
defparam \macro_inst|controller|sm_pwm|data[1] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|data[1] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[1] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[1] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[1] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[1] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[1] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[20] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[40][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan81~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [20]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~277_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [20]));
defparam \macro_inst|controller|sm_pwm|data[20] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[20] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|data[20] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[20] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[20] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[20] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[20] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[20] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[20] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[21] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan85~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[42][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [21]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~278_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [21]));
defparam \macro_inst|controller|sm_pwm|data[21] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[21] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[21] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|data[21] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[21] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[21] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[21] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[21] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[21] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[22] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmList[44][15]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan89~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [22]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y5_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~279_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [22]));
defparam \macro_inst|controller|sm_pwm|data[22] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[22] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[22] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[22] .mask = 16'h5000;
defparam \macro_inst|controller|sm_pwm|data[22] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[22] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[22] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[22] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[22] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[23] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|LessThan93~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[46][15]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [23]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~280_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [23]));
defparam \macro_inst|controller|sm_pwm|data[23] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|data[23] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[23] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|data[23] .mask = 16'h5000;
defparam \macro_inst|controller|sm_pwm|data[23] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[23] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[23] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[23] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[23] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[24] (
	.A(\macro_inst|controller|sm_pwm|LessThan1~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~216_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [24]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~217_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [24]));
defparam \macro_inst|controller|sm_pwm|data[24] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[24] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[24] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|data[24] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[24] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[24] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[24] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[24] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[24] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[25] (
	.A(\macro_inst|controller|sm_pwm|data~218_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan5~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [25]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y10_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~219_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [25]));
defparam \macro_inst|controller|sm_pwm|data[25] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|data[25] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[25] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|data[25] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[25] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[25] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[25] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[25] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[25] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[26] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|data~240_combout ),
	.C(\macro_inst|controller|sm_pwm|LessThan9~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [26]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~241_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [26]));
defparam \macro_inst|controller|sm_pwm|data[26] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[26] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[26] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[26] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[26] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[26] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[26] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[26] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[26] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[27] (
	.A(\macro_inst|controller|sm_pwm|LessThan14~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~250_combout ),
	.C(\macro_inst|controller|sm_pwm|LessThan13~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [27]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~251_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [27]));
defparam \macro_inst|controller|sm_pwm|data[27] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[27] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[27] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|data[27] .mask = 16'h2230;
defparam \macro_inst|controller|sm_pwm|data[27] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[27] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[27] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[27] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[27] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[28] (
	.A(\macro_inst|controller|sm_pwm|data~252_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan17~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [28]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y8_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~253_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [28]));
defparam \macro_inst|controller|sm_pwm|data[28] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[28] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[28] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|data[28] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[28] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[28] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[28] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[28] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[28] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[29] (
	.A(\macro_inst|controller|sm_pwm|data~254_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan21~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [29]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y10_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~255_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [29]));
defparam \macro_inst|controller|sm_pwm|data[29] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data[29] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|data[29] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[29] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[29] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[29] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[29] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[29] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[29] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[2] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[4][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan9~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~276_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [2]));
defparam \macro_inst|controller|sm_pwm|data[2] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[2] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[2] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[2] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[2] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[2] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[2] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[30] (
	.A(\macro_inst|controller|sm_pwm|data~256_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan25~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [30]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~257_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [30]));
defparam \macro_inst|controller|sm_pwm|data[30] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[30] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|data[30] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|data[30] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[30] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[30] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[30] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[30] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[30] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[31] (
	.A(\macro_inst|controller|sm_pwm|data~258_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan29~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [31]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~259_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [31]));
defparam \macro_inst|controller|sm_pwm|data[31] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[31] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[31] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[31] .mask = 16'h0504;
defparam \macro_inst|controller|sm_pwm|data[31] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[31] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[31] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[31] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[31] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[32] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|LessThan33~12_combout ),
	.D(\macro_inst|controller|sm_pwm|data~260_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [32]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~261_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [32]));
defparam \macro_inst|controller|sm_pwm|data[32] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|data[32] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[32] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|data[32] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[32] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[32] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[32] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[32] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[32] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[33] (
	.A(\macro_inst|controller|sm_pwm|data~262_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|LessThan37~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [33]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X54_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~263_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [33]));
defparam \macro_inst|controller|sm_pwm|data[33] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|data[33] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[33] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data[33] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[33] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[33] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[33] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[33] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[33] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[34] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|data~220_combout ),
	.C(\macro_inst|controller|sm_pwm|LessThan42~12_combout ),
	.D(\macro_inst|controller|sm_pwm|LessThan41~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [34]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X54_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~221_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [34]));
defparam \macro_inst|controller|sm_pwm|data[34] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[34] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data[34] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[34] .mask = 16'h3120;
defparam \macro_inst|controller|sm_pwm|data[34] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[34] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[34] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[34] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[34] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[35] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|LessThan45~12_combout ),
	.C(\macro_inst|controller|sm_pwm|data~222_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [35]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~223_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [35]));
defparam \macro_inst|controller|sm_pwm|data[35] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|data[35] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[35] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[35] .mask = 16'h0504;
defparam \macro_inst|controller|sm_pwm|data[35] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[35] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[35] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[35] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[35] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[36] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|LessThan49~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|data~224_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [36]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~225_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [36]));
defparam \macro_inst|controller|sm_pwm|data[36] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[36] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|data[36] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[36] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[36] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[36] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[36] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[36] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[36] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[37] (
	.A(\macro_inst|controller|sm_pwm|data~226_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|LessThan53~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [37]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y6_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~227_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [37]));
defparam \macro_inst|controller|sm_pwm|data[37] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[37] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[37] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[37] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[37] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[37] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[37] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[37] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[37] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[38] (
	.A(\macro_inst|controller|sm_pwm|data~228_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|LessThan57~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [38]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~229_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [38]));
defparam \macro_inst|controller|sm_pwm|data[38] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[38] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[38] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[38] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[38] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[38] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[38] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[38] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[38] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[39] (
	.A(\macro_inst|controller|sm_pwm|LessThan61~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~230_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [39]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~231_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [39]));
defparam \macro_inst|controller|sm_pwm|data[39] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[39] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|data[39] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[39] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[39] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[39] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[39] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[39] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[39] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[3] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[6][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan13~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [3]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~281_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [3]));
defparam \macro_inst|controller|sm_pwm|data[3] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[3] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[3] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|data[3] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[3] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[3] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[3] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[40] (
	.A(\macro_inst|controller|sm_pwm|LessThan65~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|data~232_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [40]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~233_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [40]));
defparam \macro_inst|controller|sm_pwm|data[40] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[40] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|data[40] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[40] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[40] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[40] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[40] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[40] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[40] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[41] (
	.A(\macro_inst|controller|sm_pwm|LessThan69~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|LessThan70~12_combout ),
	.D(\macro_inst|controller|sm_pwm|data~234_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [41]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~235_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [41]));
defparam \macro_inst|controller|sm_pwm|data[41] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[41] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data[41] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[41] .mask = 16'h00E2;
defparam \macro_inst|controller|sm_pwm|data[41] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[41] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[41] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[41] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[41] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[42] (
	.A(\macro_inst|controller|sm_pwm|data~236_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan73~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [42]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~237_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [42]));
defparam \macro_inst|controller|sm_pwm|data[42] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[42] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[42] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|data[42] .mask = 16'h0504;
defparam \macro_inst|controller|sm_pwm|data[42] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[42] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[42] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[42] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[42] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[43] (
	.A(\macro_inst|controller|sm_pwm|data~238_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan77~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [43]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y5_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~239_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [43]));
defparam \macro_inst|controller|sm_pwm|data[43] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[43] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|data[43] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|data[43] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[43] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[43] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[43] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[43] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[43] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[44] (
	.A(\macro_inst|controller|sm_pwm|data~242_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan81~12_combout ),
	.C(\macro_inst|controller|sm_pwm|LessThan82~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [44]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~243_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [44]));
defparam \macro_inst|controller|sm_pwm|data[44] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[44] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|data[44] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|data[44] .mask = 16'h5044;
defparam \macro_inst|controller|sm_pwm|data[44] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[44] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[44] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[44] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[44] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[45] (
	.A(\macro_inst|controller|sm_pwm|data~244_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan85~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [45]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~245_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [45]));
defparam \macro_inst|controller|sm_pwm|data[45] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[45] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[45] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[45] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[45] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[45] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[45] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[45] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[45] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[46] (
	.A(\macro_inst|controller|sm_pwm|data~246_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan89~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [46]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y5_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~247_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [46]));
defparam \macro_inst|controller|sm_pwm|data[46] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[46] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[46] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[46] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[46] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[46] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[46] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[46] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[46] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[47] (
	.A(\macro_inst|controller|sm_pwm|data~248_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|LessThan93~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [47]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~249_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [47]));
defparam \macro_inst|controller|sm_pwm|data[47] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|data[47] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[47] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[47] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[47] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[47] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[47] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[47] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[47] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[48] (
	.A(\macro_inst|controller|sm_pwm|LessThan2~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~168_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [48]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~169_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [48]));
defparam \macro_inst|controller|sm_pwm|data[48] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[48] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[48] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[48] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[48] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[48] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[48] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[48] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[48] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[49] (
	.A(\macro_inst|controller|sm_pwm|data~170_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan6~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [49]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y10_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~171_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [49]));
defparam \macro_inst|controller|sm_pwm|data[49] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|data[49] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[49] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[49] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[49] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[49] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[49] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[49] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[49] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[8][15]~q ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|LessThan17~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [4]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~282_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [4]));
defparam \macro_inst|controller|sm_pwm|data[4] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[4] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[4] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|data[4] .mask = 16'h00A0;
defparam \macro_inst|controller|sm_pwm|data[4] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[4] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[4] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[50] (
	.A(\macro_inst|controller|sm_pwm|LessThan10~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|data~192_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [50]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~193_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [50]));
defparam \macro_inst|controller|sm_pwm|data[50] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[50] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[50] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|data[50] .mask = 16'h000E;
defparam \macro_inst|controller|sm_pwm|data[50] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[50] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[50] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[50] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[50] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[51] (
	.A(\macro_inst|controller|sm_pwm|LessThan14~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|data~202_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [51]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~203_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [51]));
defparam \macro_inst|controller|sm_pwm|data[51] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[51] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[51] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|data[51] .mask = 16'h000E;
defparam \macro_inst|controller|sm_pwm|data[51] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[51] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[51] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[51] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[51] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[52] (
	.A(\macro_inst|controller|sm_pwm|LessThan18~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~204_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|LessThan17~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [52]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y8_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~205_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [52]));
defparam \macro_inst|controller|sm_pwm|data[52] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[52] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[52] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|data[52] .mask = 16'h3202;
defparam \macro_inst|controller|sm_pwm|data[52] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[52] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[52] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[52] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[52] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[53] (
	.A(\macro_inst|controller|sm_pwm|LessThan22~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~206_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [53]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y10_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~207_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [53]));
defparam \macro_inst|controller|sm_pwm|data[53] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data[53] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|data[53] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[53] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[53] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[53] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[53] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[53] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[53] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[54] (
	.A(\macro_inst|controller|sm_pwm|data~208_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan26~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [54]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~209_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [54]));
defparam \macro_inst|controller|sm_pwm|data[54] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[54] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|data[54] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|data[54] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[54] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[54] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[54] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[54] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[54] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[55] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|LessThan30~12_combout ),
	.C(\macro_inst|controller|sm_pwm|data~210_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [55]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~211_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [55]));
defparam \macro_inst|controller|sm_pwm|data[55] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[55] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[55] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[55] .mask = 16'h000E;
defparam \macro_inst|controller|sm_pwm|data[55] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[55] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[55] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[55] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[55] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[56] (
	.A(\macro_inst|controller|sm_pwm|data~212_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|LessThan34~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [56]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~213_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [56]));
defparam \macro_inst|controller|sm_pwm|data[56] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|data[56] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[56] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|data[56] .mask = 16'h0504;
defparam \macro_inst|controller|sm_pwm|data[56] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[56] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[56] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[56] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[56] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[57] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|LessThan38~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|data~214_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [57]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X54_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~215_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [57]));
defparam \macro_inst|controller|sm_pwm|data[57] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|data[57] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[57] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|data[57] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[57] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[57] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[57] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[57] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[57] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[58] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|data~172_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|LessThan42~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [58]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X54_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~173_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [58]));
defparam \macro_inst|controller|sm_pwm|data[58] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[58] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data[58] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|data[58] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[58] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[58] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[58] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[58] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[58] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[59] (
	.A(\macro_inst|controller|sm_pwm|LessThan46~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|data~174_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [59]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~175_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [59]));
defparam \macro_inst|controller|sm_pwm|data[59] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|data[59] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[59] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|data[59] .mask = 16'h0302;
defparam \macro_inst|controller|sm_pwm|data[59] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[59] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[59] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[59] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[59] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[5] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan21~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[10][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [5]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y10_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~283_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [5]));
defparam \macro_inst|controller|sm_pwm|data[5] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data[5] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|data[5] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[5] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[60] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|LessThan50~12_combout ),
	.C(\macro_inst|controller|sm_pwm|data~176_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [60]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~177_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [60]));
defparam \macro_inst|controller|sm_pwm|data[60] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[60] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|data[60] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|data[60] .mask = 16'h000E;
defparam \macro_inst|controller|sm_pwm|data[60] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[60] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[60] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[60] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[60] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[61] (
	.A(\macro_inst|controller|sm_pwm|LessThan53~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|LessThan54~12_combout ),
	.D(\macro_inst|controller|sm_pwm|data~178_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [61]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y6_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~179_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [61]));
defparam \macro_inst|controller|sm_pwm|data[61] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[61] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[61] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|data[61] .mask = 16'h00B8;
defparam \macro_inst|controller|sm_pwm|data[61] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[61] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[61] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[61] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[61] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[62] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|data~180_combout ),
	.C(\macro_inst|controller|sm_pwm|LessThan58~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [62]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~181_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [62]));
defparam \macro_inst|controller|sm_pwm|data[62] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[62] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[62] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[62] .mask = 16'h1110;
defparam \macro_inst|controller|sm_pwm|data[62] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[62] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[62] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[62] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[62] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[63] (
	.A(\macro_inst|controller|sm_pwm|LessThan62~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~182_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [63]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~183_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [63]));
defparam \macro_inst|controller|sm_pwm|data[63] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[63] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|data[63] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[63] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[63] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[63] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[63] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[63] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[63] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[64] (
	.A(\macro_inst|controller|sm_pwm|data~184_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan66~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [64]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~185_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [64]));
defparam \macro_inst|controller|sm_pwm|data[64] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[64] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|data[64] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data[64] .mask = 16'h0504;
defparam \macro_inst|controller|sm_pwm|data[64] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[64] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[64] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[64] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[64] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[65] (
	.A(\macro_inst|controller|sm_pwm|data~186_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|LessThan70~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [65]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~187_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [65]));
defparam \macro_inst|controller|sm_pwm|data[65] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[65] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data[65] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[65] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[65] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[65] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[65] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[65] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[65] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[66] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|LessThan74~12_combout ),
	.C(\macro_inst|controller|sm_pwm|data~188_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [66]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~189_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [66]));
defparam \macro_inst|controller|sm_pwm|data[66] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[66] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data[66] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[66] .mask = 16'h0504;
defparam \macro_inst|controller|sm_pwm|data[66] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[66] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[66] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[66] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[66] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[67] (
	.A(\macro_inst|controller|sm_pwm|LessThan78~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~190_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [67]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y5_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~191_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [67]));
defparam \macro_inst|controller|sm_pwm|data[67] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[67] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|data[67] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|data[67] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[67] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[67] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[67] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[67] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[67] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[68] (
	.A(\macro_inst|controller|sm_pwm|LessThan82~12_combout ),
	.B(\macro_inst|controller|sm_pwm|data~194_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [68]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~195_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [68]));
defparam \macro_inst|controller|sm_pwm|data[68] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[68] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|data[68] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data[68] .mask = 16'h0032;
defparam \macro_inst|controller|sm_pwm|data[68] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[68] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[68] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[68] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[68] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[69] (
	.A(\macro_inst|controller|sm_pwm|data~196_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan86~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [69]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~197_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [69]));
defparam \macro_inst|controller|sm_pwm|data[69] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[69] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[69] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|data[69] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[69] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[69] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[69] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[69] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[69] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[6] (
	.A(\macro_inst|controller|sm_pwm|LessThan25~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[12][15]~q ),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [6]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~284_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [6]));
defparam \macro_inst|controller|sm_pwm|data[6] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[6] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|data[6] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[6] .mask = 16'h0088;
defparam \macro_inst|controller|sm_pwm|data[6] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[6] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[70] (
	.A(\macro_inst|controller|sm_pwm|data~198_combout ),
	.B(\macro_inst|controller|sm_pwm|LessThan90~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [70]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y5_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~199_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [70]));
defparam \macro_inst|controller|sm_pwm|data[70] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[70] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[70] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[70] .mask = 16'h0054;
defparam \macro_inst|controller|sm_pwm|data[70] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[70] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[70] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[70] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[70] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[71] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|data~200_combout ),
	.D(\macro_inst|controller|sm_pwm|LessThan94~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [71]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~201_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [71]));
defparam \macro_inst|controller|sm_pwm|data[71] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|data[71] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[71] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data[71] .mask = 16'h0504;
defparam \macro_inst|controller|sm_pwm|data[71] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[71] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[71] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[71] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[71] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[72] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[0][7]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan2~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [72]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~144_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [72]));
defparam \macro_inst|controller|sm_pwm|data[72] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[72] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[72] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[72] .mask = 16'h0030;
defparam \macro_inst|controller|sm_pwm|data[72] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[72] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[72] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[72] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[72] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[73] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan6~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[2][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [73]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y10_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~145_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [73]));
defparam \macro_inst|controller|sm_pwm|data[73] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|data[73] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[73] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[73] .mask = 16'h000C;
defparam \macro_inst|controller|sm_pwm|data[73] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[73] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[73] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[73] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[73] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[74] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[4][7]~q ),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|LessThan10~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [74]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y12_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~156_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [74]));
defparam \macro_inst|controller|sm_pwm|data[74] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[74] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[74] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[74] .mask = 16'h0300;
defparam \macro_inst|controller|sm_pwm|data[74] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[74] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[74] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[74] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[74] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[75] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[6][7]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan14~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [75]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~161_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [75]));
defparam \macro_inst|controller|sm_pwm|data[75] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[75] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[75] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|data[75] .mask = 16'h0030;
defparam \macro_inst|controller|sm_pwm|data[75] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[75] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[75] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[75] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[75] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[76] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[8][7]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan18~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [76]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y8_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~162_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [76]));
defparam \macro_inst|controller|sm_pwm|data[76] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[76] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[76] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|data[76] .mask = 16'h0030;
defparam \macro_inst|controller|sm_pwm|data[76] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[76] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[76] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[76] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[76] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[77] (
	.A(\macro_inst|controller|sm_pwm|LessThan22~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[10][7]~q ),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [77]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y10_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~163_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [77]));
defparam \macro_inst|controller|sm_pwm|data[77] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data[77] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|data[77] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|data[77] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|data[77] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[77] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[77] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[77] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[77] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[78] (
	.A(\macro_inst|controller|sm_pwm|pwmList[12][7]~q ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|LessThan26~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [78]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~164_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [78]));
defparam \macro_inst|controller|sm_pwm|data[78] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[78] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|data[78] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data[78] .mask = 16'h0050;
defparam \macro_inst|controller|sm_pwm|data[78] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[78] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[78] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[78] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[78] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[79] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[14][7]~q ),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|LessThan30~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [79]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~165_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [79]));
defparam \macro_inst|controller|sm_pwm|data[79] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[79] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[79] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|data[79] .mask = 16'h0300;
defparam \macro_inst|controller|sm_pwm|data[79] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[79] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[79] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[79] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[79] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[7] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|LessThan29~12_combout ),
	.C(vcc),
	.D(\macro_inst|controller|sm_pwm|pwmList[14][15]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [7]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~285_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [7]));
defparam \macro_inst|controller|sm_pwm|data[7] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[7] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[7] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|data[7] .mask = 16'h4400;
defparam \macro_inst|controller|sm_pwm|data[7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[80] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan34~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|pwmList[16][7]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [80]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~166_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [80]));
defparam \macro_inst|controller|sm_pwm|data[80] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|data[80] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[80] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[80] .mask = 16'h000C;
defparam \macro_inst|controller|sm_pwm|data[80] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[80] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[80] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[80] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[80] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[81] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[18][7]~q ),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|LessThan38~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [81]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X54_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~167_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [81]));
defparam \macro_inst|controller|sm_pwm|data[81] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|data[81] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[81] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|data[81] .mask = 16'h0300;
defparam \macro_inst|controller|sm_pwm|data[81] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[81] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[81] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[81] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[81] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[82] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|pwmList[20][7]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan42~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [82]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X54_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~146_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [82]));
defparam \macro_inst|controller|sm_pwm|data[82] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[82] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data[82] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[82] .mask = 16'h0300;
defparam \macro_inst|controller|sm_pwm|data[82] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[82] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[82] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[82] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[82] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[83] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmList[22][7]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan46~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [83]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~147_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [83]));
defparam \macro_inst|controller|sm_pwm|data[83] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|data[83] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[83] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data[83] .mask = 16'h0500;
defparam \macro_inst|controller|sm_pwm|data[83] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[83] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[83] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[83] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[83] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[84] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[24][7]~q ),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|LessThan50~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [84]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~148_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [84]));
defparam \macro_inst|controller|sm_pwm|data[84] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[84] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|data[84] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data[84] .mask = 16'h0300;
defparam \macro_inst|controller|sm_pwm|data[84] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[84] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[84] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[84] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[84] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[85] (
	.A(\macro_inst|controller|sm_pwm|pwmList[26][7]~q ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|LessThan54~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [85]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y6_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~149_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [85]));
defparam \macro_inst|controller|sm_pwm|data[85] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[85] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[85] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[85] .mask = 16'h0050;
defparam \macro_inst|controller|sm_pwm|data[85] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[85] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[85] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[85] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[85] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[86] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan58~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[28][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [86]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~150_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [86]));
defparam \macro_inst|controller|sm_pwm|data[86] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[86] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[86] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|data[86] .mask = 16'h000C;
defparam \macro_inst|controller|sm_pwm|data[86] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[86] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[86] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[86] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[86] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[87] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|pwmList[30][7]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan62~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [87]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X56_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~151_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [87]));
defparam \macro_inst|controller|sm_pwm|data[87] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[87] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|data[87] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|data[87] .mask = 16'h0300;
defparam \macro_inst|controller|sm_pwm|data[87] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[87] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[87] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[87] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[87] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[88] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[32][7]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan66~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [88]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~152_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [88]));
defparam \macro_inst|controller|sm_pwm|data[88] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[88] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|data[88] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|data[88] .mask = 16'h0030;
defparam \macro_inst|controller|sm_pwm|data[88] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[88] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[88] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[88] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[88] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[89] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[34][7]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan70~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [89]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~153_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [89]));
defparam \macro_inst|controller|sm_pwm|data[89] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data[89] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data[89] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[89] .mask = 16'h0030;
defparam \macro_inst|controller|sm_pwm|data[89] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[89] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[89] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[89] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[89] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[8] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|LessThan33~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[16][15]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [8]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~286_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [8]));
defparam \macro_inst|controller|sm_pwm|data[8] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|data[8] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[8] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data[8] .mask = 16'h5000;
defparam \macro_inst|controller|sm_pwm|data[8] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[8] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[8] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[90] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan74~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[36][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [90]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X58_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~154_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [90]));
defparam \macro_inst|controller|sm_pwm|data[90] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[90] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data[90] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|data[90] .mask = 16'h000C;
defparam \macro_inst|controller|sm_pwm|data[90] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[90] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[90] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[90] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[90] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[91] (
	.A(\macro_inst|controller|sm_pwm|LessThan78~12_combout ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmList[38][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [91]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y5_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~155_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [91]));
defparam \macro_inst|controller|sm_pwm|data[91] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[91] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|data[91] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|data[91] .mask = 16'h000A;
defparam \macro_inst|controller|sm_pwm|data[91] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[91] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[91] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[91] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[91] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[92] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[40][7]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan82~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [92]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y9_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~157_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [92]));
defparam \macro_inst|controller|sm_pwm|data[92] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[92] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|data[92] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[92] .mask = 16'h0030;
defparam \macro_inst|controller|sm_pwm|data[92] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[92] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[92] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[92] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[92] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[93] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan86~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[42][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [93]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X62_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~158_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [93]));
defparam \macro_inst|controller|sm_pwm|data[93] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[93] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data[93] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|data[93] .mask = 16'h000C;
defparam \macro_inst|controller|sm_pwm|data[93] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[93] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[93] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[93] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[93] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[94] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan90~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[44][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [94]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y5_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~159_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [94]));
defparam \macro_inst|controller|sm_pwm|data[94] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data[94] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[94] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data[94] .mask = 16'h000C;
defparam \macro_inst|controller|sm_pwm|data[94] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[94] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[94] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[94] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[94] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[95] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmList[46][7]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan94~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [95]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y1_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~160_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [95]));
defparam \macro_inst|controller|sm_pwm|data[95] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|data[95] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[95] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|data[95] .mask = 16'h0500;
defparam \macro_inst|controller|sm_pwm|data[95] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[95] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[95] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[95] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[95] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[96] (
	.A(\macro_inst|controller|sm_pwm|LessThan3~12_combout ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|pwmList[1][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [96]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~120_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [96]));
defparam \macro_inst|controller|sm_pwm|data[96] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data[96] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[96] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data[96] .mask = 16'h00A0;
defparam \macro_inst|controller|sm_pwm|data[96] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[96] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[96] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[96] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[96] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[97] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(\macro_inst|controller|sm_pwm|pwmList[3][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan7~12_combout ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [97]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X57_Y7_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~121_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [97]));
defparam \macro_inst|controller|sm_pwm|data[97] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data[97] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data[97] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|data[97] .mask = 16'h4040;
defparam \macro_inst|controller|sm_pwm|data[97] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[97] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[97] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[97] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[97] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[98] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan11~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[5][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [98]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X61_Y11_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~132_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [98]));
defparam \macro_inst|controller|sm_pwm|data[98] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data[98] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data[98] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data[98] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[98] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[98] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[98] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[98] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[98] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[99] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|LessThan15~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[7][15]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [99]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X60_Y6_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~137_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [99]));
defparam \macro_inst|controller|sm_pwm|data[99] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data[99] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|data[99] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|data[99] .mask = 16'h5000;
defparam \macro_inst|controller|sm_pwm|data[99] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[99] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[99] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[99] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[99] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data[9] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|LessThan37~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[18][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|data [9]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X54_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~287_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|data [9]));
defparam \macro_inst|controller|sm_pwm|data[9] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|data[9] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data[9] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|data[9] .mask = 16'h00C0;
defparam \macro_inst|controller|sm_pwm|data[9] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[9] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data[9] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~100 (
	.A(\macro_inst|controller|sm_pwm|LessThan88~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[43][15]~q ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmList[43][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~100_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~100 .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data~100 .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data~100 .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|data~100 .mask = 16'h5CFC;
defparam \macro_inst|controller|sm_pwm|data~100 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~100 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~100 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~100 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~100 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~102 (
	.A(\macro_inst|controller|sm_pwm|pwmList[45][7]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmList[45][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan92~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~102_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~102 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data~102 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data~102 .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|data~102 .mask = 16'h5FCC;
defparam \macro_inst|controller|sm_pwm|data~102 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~102 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~102 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~102 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~102 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~106 (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|LessThan16~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[7][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmList[7][15]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~106_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~106 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data~106 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|data~106 .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data~106 .mask = 16'h7F2A;
defparam \macro_inst|controller|sm_pwm|data~106 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~106 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~106 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~106 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~106 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~108 (
	.A(\macro_inst|controller|sm_pwm|pwmList[9][7]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan20~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmList[9][15]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~108_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~108 .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data~108 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data~108 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|data~108 .mask = 16'h7F70;
defparam \macro_inst|controller|sm_pwm|data~108 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~108 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~108 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~108 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~108 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~112 (
	.A(\macro_inst|controller|sm_pwm|pwmList[13][15]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmList[13][7]~q ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|LessThan28~12_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~112_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~112 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data~112 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data~112 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data~112 .mask = 16'h3AFA;
defparam \macro_inst|controller|sm_pwm|data~112 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~112 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~112 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~112 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~112 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~116 (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[17][7]~q ),
	.C(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.D(\macro_inst|controller|sm_pwm|pwmList[17][15]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~116_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~116 .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|data~116 .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data~116 .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data~116 .mask = 16'hF7F2;
defparam \macro_inst|controller|sm_pwm|data~116 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~116 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~116 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~116 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~116 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~118 (
	.A(\macro_inst|controller|sm_pwm|LessThan40~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|pwmList[19][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmList[19][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~118_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~118 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data~118 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data~118 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|data~118 .mask = 16'h74FC;
defparam \macro_inst|controller|sm_pwm|data~118 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~118 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~118 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~118 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~118 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~168 (
	.A(\macro_inst|controller|sm_pwm|pwmList[0][15]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|LessThan1~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[0][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~168_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~168 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data~168 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data~168 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|data~168 .mask = 16'h8CBF;
defparam \macro_inst|controller|sm_pwm|data~168 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~168 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~168 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~168 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~168 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~170 (
	.A(\macro_inst|controller|sm_pwm|LessThan5~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|pwmList[2][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmList[2][15]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~170_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~170 .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|data~170 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data~170 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|data~170 .mask = 16'hCF47;
defparam \macro_inst|controller|sm_pwm|data~170 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~170 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~170 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~170 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~170 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~172 (
	.A(\macro_inst|controller|sm_pwm|pwmList[20][15]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|pwmList[20][7]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan41~12_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~172_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~172 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data~172 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data~172 .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data~172 .mask = 16'h8BCF;
defparam \macro_inst|controller|sm_pwm|data~172 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~172 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~172 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~172 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~172 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~176 (
	.A(\macro_inst|controller|sm_pwm|LessThan49~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[24][15]~q ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmList[24][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~176_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~176 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data~176 .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|data~176 .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data~176 .mask = 16'hD0DF;
defparam \macro_inst|controller|sm_pwm|data~176 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~176 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~176 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~176 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~176 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~182 (
	.A(\macro_inst|controller|sm_pwm|pwmList[30][15]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|LessThan61~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[30][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~182_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~182 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data~182 .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|data~182 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|data~182 .mask = 16'h8CBF;
defparam \macro_inst|controller|sm_pwm|data~182 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~182 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~182 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~182 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~182 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~186 (
	.A(\macro_inst|controller|sm_pwm|LessThan69~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|pwmList[34][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmList[34][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~186_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~186 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data~186 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data~186 .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data~186 .mask = 16'hC4F7;
defparam \macro_inst|controller|sm_pwm|data~186 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~186 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~186 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~186 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~186 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~190 (
	.A(\macro_inst|controller|sm_pwm|pwmList[38][7]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|LessThan77~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[38][15]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~190_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~190 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data~190 .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|data~190 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|data~190 .mask = 16'hDD1D;
defparam \macro_inst|controller|sm_pwm|data~190 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~190 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~190 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~190 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~190 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~192 (
	.A(\macro_inst|controller|sm_pwm|pwmList[4][7]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmList[4][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan9~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~192_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~192 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data~192 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data~192 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|data~192 .mask = 16'hCF55;
defparam \macro_inst|controller|sm_pwm|data~192 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~192 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~192 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~192 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~192 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~194 (
	.A(\macro_inst|controller|sm_pwm|pwmList[40][7]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan81~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmList[40][15]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~194_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~194 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data~194 .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|data~194 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|data~194 .mask = 16'hF535;
defparam \macro_inst|controller|sm_pwm|data~194 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~194 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~194 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~194 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~194 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~200 (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|LessThan93~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[46][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmList[46][15]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~200_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~200 .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|data~200 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data~200 .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|data~200 .mask = 16'hAF27;
defparam \macro_inst|controller|sm_pwm|data~200 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~200 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~200 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~200 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~200 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~214 (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|LessThan37~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[18][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmList[18][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~214_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~214 .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|data~214 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data~214 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|data~214 .mask = 16'hA2F7;
defparam \macro_inst|controller|sm_pwm|data~214 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~214 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~214 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~214 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~214 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~218 (
	.A(\macro_inst|controller|sm_pwm|pwmList[2][7]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmList[2][15]~q ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|LessThan6~12_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~218_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~218 .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|data~218 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data~218 .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data~218 .mask = 16'h5CFC;
defparam \macro_inst|controller|sm_pwm|data~218 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~218 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~218 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~218 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~218 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~220 (
	.A(\macro_inst|controller|sm_pwm|pwmList[20][7]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|pwmList[20][15]~q ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~220_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~220 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data~220 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data~220 .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|data~220 .mask = 16'hDDFC;
defparam \macro_inst|controller|sm_pwm|data~220 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~220 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~220 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~220 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~220 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~224 (
	.A(\macro_inst|controller|sm_pwm|LessThan50~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[24][7]~q ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmList[24][15]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~224_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~224 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data~224 .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|data~224 .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|data~224 .mask = 16'h7F70;
defparam \macro_inst|controller|sm_pwm|data~224 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~224 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~224 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~224 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~224 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~226 (
	.A(\macro_inst|controller|sm_pwm|pwmList[26][7]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|LessThan54~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[26][15]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~226_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~226 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data~226 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data~226 .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data~226 .mask = 16'h7F4C;
defparam \macro_inst|controller|sm_pwm|data~226 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~226 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~226 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~226 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~226 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~234 (
	.A(\macro_inst|controller|sm_pwm|pwmList[34][15]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmList[34][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~234_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~234 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data~234 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data~234 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|data~234 .mask = 16'hCEFE;
defparam \macro_inst|controller|sm_pwm|data~234 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~234 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~234 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~234 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~234 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~248 (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|LessThan94~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[46][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmList[46][15]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~248_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~248 .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|data~248 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data~248 .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|data~248 .mask = 16'h7F2A;
defparam \macro_inst|controller|sm_pwm|data~248 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~248 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~248 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~248 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~248 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~26 (
	.A(\macro_inst|controller|sm_pwm|LessThan7~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[3][15]~q ),
	.C(\macro_inst|controller|sm_pwm|pwmList[3][7]~q ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~26_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~26 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data~26 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data~26 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data~26 .mask = 16'hDD0F;
defparam \macro_inst|controller|sm_pwm|data~26 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~26 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~26 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~26 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~26 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~28 (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[21][15]~q ),
	.C(\macro_inst|controller|sm_pwm|pwmList[21][7]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan43~12_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~28_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~28 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data~28 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|data~28 .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data~28 .mask = 16'h8DAF;
defparam \macro_inst|controller|sm_pwm|data~28 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~28 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~28 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~28 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~28 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~32 (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[25][15]~q ),
	.C(\macro_inst|controller|sm_pwm|pwmList[25][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~32_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~32 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data~32 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data~32 .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data~32 .mask = 16'hFF8D;
defparam \macro_inst|controller|sm_pwm|data~32 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~32 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~32 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~32 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~32 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~34 (
	.A(\macro_inst|controller|sm_pwm|pwmList[27][15]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmList[27][7]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan55~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~34_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~34 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data~34 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data~34 .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data~34 .mask = 16'hAF33;
defparam \macro_inst|controller|sm_pwm|data~34 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~34 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~34 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~34 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~34 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~36 (
	.A(\macro_inst|controller|sm_pwm|pwmList[29][7]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmList[29][15]~q ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|LessThan59~12_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~36_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~36 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data~36 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data~36 .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|data~36 .mask = 16'hC5F5;
defparam \macro_inst|controller|sm_pwm|data~36 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~36 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~36 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~36 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~36 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~44 (
	.A(\macro_inst|controller|sm_pwm|pwmList[37][15]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan75~12_combout ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmList[37][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~44_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~44 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data~44 .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data~44 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data~44 .mask = 16'hB0BF;
defparam \macro_inst|controller|sm_pwm|data~44 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~44 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~44 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~44 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~44 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~46 (
	.A(\macro_inst|controller|sm_pwm|LessThan79~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|pwmList[39][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmList[39][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~46_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~46 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data~46 .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|data~46 .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|data~46 .mask = 16'hC4F7;
defparam \macro_inst|controller|sm_pwm|data~46 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~46 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~46 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~46 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~46 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~48 (
	.A(\macro_inst|controller|sm_pwm|pwmList[5][15]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmList[5][7]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan11~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~48_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~48 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data~48 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data~48 .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|data~48 .mask = 16'hAF33;
defparam \macro_inst|controller|sm_pwm|data~48 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~48 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~48 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~48 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~48 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~50 (
	.A(\macro_inst|controller|sm_pwm|pwmList[41][7]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmList[41][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan83~12_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~50_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~50 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data~50 .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|data~50 .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data~50 .mask = 16'hCF55;
defparam \macro_inst|controller|sm_pwm|data~50 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~50 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~50 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~50 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~50 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~52 (
	.A(\macro_inst|controller|sm_pwm|pwmList[43][7]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan87~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[43][15]~q ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~52_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~52 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data~52 .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|data~52 .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|data~52 .mask = 16'hF355;
defparam \macro_inst|controller|sm_pwm|data~52 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~52 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~52 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~52 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~52 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~54 (
	.A(\macro_inst|controller|sm_pwm|LessThan91~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|pwmList[45][15]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmList[45][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~54_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~54 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data~54 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data~54 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data~54 .mask = 16'hC4F7;
defparam \macro_inst|controller|sm_pwm|data~54 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~54 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~54 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~54 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~54 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~60 (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|LessThan19~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[9][7]~q ),
	.D(\macro_inst|controller|sm_pwm|pwmList[9][15]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~60_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~60 .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|data~60 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data~60 .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data~60 .mask = 16'hAF27;
defparam \macro_inst|controller|sm_pwm|data~60 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~60 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~60 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~60 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~60 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~64 (
	.A(\macro_inst|controller|sm_pwm|pwmList[13][15]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmList[13][7]~q ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~64_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~64 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data~64 .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|data~64 .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data~64 .mask = 16'hFFA3;
defparam \macro_inst|controller|sm_pwm|data~64 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~64 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~64 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~64 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~64 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~66 (
	.A(\macro_inst|controller|sm_pwm|pwmList[15][15]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|LessThan31~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[15][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~66_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~66 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data~66 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data~66 .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data~66 .mask = 16'h8CBF;
defparam \macro_inst|controller|sm_pwm|data~66 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~66 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~66 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~66 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~66 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~68 (
	.A(\macro_inst|controller|sm_pwm|LessThan35~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[17][7]~q ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|pwmList[17][15]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~68_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~68 .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|data~68 .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|data~68 .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|data~68 .mask = 16'hF353;
defparam \macro_inst|controller|sm_pwm|data~68 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~68 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~68 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~68 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~68 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~70 (
	.A(\macro_inst|controller|sm_pwm|pwmList[19][7]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan39~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[19][15]~q ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~70_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~70 .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|data~70 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data~70 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|data~70 .mask = 16'hF355;
defparam \macro_inst|controller|sm_pwm|data~70 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~70 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~70 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~70 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~70 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~74 (
	.A(\macro_inst|controller|sm_pwm|pwmList[3][7]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\macro_inst|controller|sm_pwm|pwmList[3][15]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan8~12_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~74_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~74 .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|data~74 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|data~74 .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|data~74 .mask = 16'h74FC;
defparam \macro_inst|controller|sm_pwm|data~74 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~74 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~74 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~74 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~74 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~78 (
	.A(\macro_inst|controller|sm_pwm|pwmList[23][15]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan48~12_combout ),
	.C(\macro_inst|controller|sm_pwm|pwmList[23][7]~q ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~78_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~78 .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|data~78 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|data~78 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data~78 .mask = 16'h3FAA;
defparam \macro_inst|controller|sm_pwm|data~78 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~78 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~78 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~78 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~78 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~80 (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[25][15]~q ),
	.C(\macro_inst|controller|sm_pwm|pwmList[25][7]~q ),
	.D(\macro_inst|controller|sm_pwm|LessThan52~12_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~80_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~80 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|data~80 .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|data~80 .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|data~80 .mask = 16'h4EEE;
defparam \macro_inst|controller|sm_pwm|data~80 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~80 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~80 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~80 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~80 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~90 (
	.A(\macro_inst|controller|sm_pwm|pwmList[35][7]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmList[35][15]~q ),
	.C(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.D(\macro_inst|controller|sm_pwm|LessThan72~12_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~90_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~90 .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|data~90 .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|data~90 .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|data~90 .mask = 16'h5CFC;
defparam \macro_inst|controller|sm_pwm|data~90 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~90 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~90 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~90 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~90 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~96 (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[5][15]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan12~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[5][7]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~96_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~96 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data~96 .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|data~96 .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|data~96 .mask = 16'h4EEE;
defparam \macro_inst|controller|sm_pwm|data~96 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~96 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~96 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~96 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~96 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|data~98 (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[41][7]~q ),
	.C(\macro_inst|controller|sm_pwm|LessThan84~12_combout ),
	.D(\macro_inst|controller|sm_pwm|pwmList[41][15]~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|data~98_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|data~98 .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|data~98 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|data~98 .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|data~98 .mask = 16'h7F2A;
defparam \macro_inst|controller|sm_pwm|data~98 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~98 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~98 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~98 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|data~98 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|motor_flags[0] (
	.A(\macro_inst|controller|sm_pwm|motor_flags[0]~3_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags[0]~6_combout ),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X59_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|motor_flags[0]~7_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|motor_flags [0]));
defparam \macro_inst|controller|sm_pwm|motor_flags[0] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|motor_flags[0] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|motor_flags[0] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|motor_flags[0] .mask = 16'h70F8;
defparam \macro_inst|controller|sm_pwm|motor_flags[0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|motor_flags[0] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|motor_flags[0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|motor_flags[0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|motor_flags[0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|motor_flags[0]~3 (
	.A(\macro_inst|controller|sm_pwm|motor_flags[0]~1_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags[0]~0_combout ),
	.C(\macro_inst|controller|sm_pwm|LessThan0~0_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags[0]~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|motor_flags[0]~3_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~3 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~3 .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~3 .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~3 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~3 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~3 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~3 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~3 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~3 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|motor_flags[0]~6 (
	.A(\macro_inst|controller|sm_pwm|Decoder0~5_combout ),
	.B(\macro_inst|controller|sm_pwm|Equal0~1_combout ),
	.C(\macro_inst|controller|sm_pwm|Equal0~0_combout ),
	.D(\macro_inst|controller|sm_pwm|motor_flags[0]~5_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|motor_flags[0]~6_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~6 .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~6 .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~6 .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~6 .mask = 16'h8000;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~6 .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~6 .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~6 .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~6 .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|motor_flags[0]~6 .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmCnt[0] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|pwmUpdateTrigger~q_X59_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Add0~0_combout ),
	.Cout(\macro_inst|controller|sm_pwm|Add0~1 ),
	.Q(\macro_inst|controller|sm_pwm|pwmCnt [0]));
defparam \macro_inst|controller|sm_pwm|pwmCnt[0] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmCnt[0] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmCnt[0] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmCnt[0] .mask = 16'h33CC;
defparam \macro_inst|controller|sm_pwm|pwmCnt[0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[0] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmCnt[1] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|Add0~1 ),
	.Qin(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|pwmUpdateTrigger~q_X59_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Add0~2_combout ),
	.Cout(\macro_inst|controller|sm_pwm|Add0~3 ),
	.Q(\macro_inst|controller|sm_pwm|pwmCnt [1]));
defparam \macro_inst|controller|sm_pwm|pwmCnt[1] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmCnt[1] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmCnt[1] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmCnt[1] .mask = 16'h3C3F;
defparam \macro_inst|controller|sm_pwm|pwmCnt[1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmCnt[1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[1] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmCnt[2] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|Add0~3 ),
	.Qin(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|pwmUpdateTrigger~q_X59_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Add0~4_combout ),
	.Cout(\macro_inst|controller|sm_pwm|Add0~5 ),
	.Q(\macro_inst|controller|sm_pwm|pwmCnt [2]));
defparam \macro_inst|controller|sm_pwm|pwmCnt[2] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmCnt[2] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmCnt[2] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmCnt[2] .mask = 16'hC30C;
defparam \macro_inst|controller|sm_pwm|pwmCnt[2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmCnt[2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[2] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmCnt[3] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|Add0~5 ),
	.Qin(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|pwmUpdateTrigger~q_X59_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Add0~6_combout ),
	.Cout(\macro_inst|controller|sm_pwm|Add0~7 ),
	.Q(\macro_inst|controller|sm_pwm|pwmCnt [3]));
defparam \macro_inst|controller|sm_pwm|pwmCnt[3] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmCnt[3] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmCnt[3] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmCnt[3] .mask = 16'h3C3F;
defparam \macro_inst|controller|sm_pwm|pwmCnt[3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmCnt[3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[3] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmCnt[4] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|Add0~7 ),
	.Qin(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|pwmUpdateTrigger~q_X59_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Add0~8_combout ),
	.Cout(\macro_inst|controller|sm_pwm|Add0~9 ),
	.Q(\macro_inst|controller|sm_pwm|pwmCnt [4]));
defparam \macro_inst|controller|sm_pwm|pwmCnt[4] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmCnt[4] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmCnt[4] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmCnt[4] .mask = 16'hC30C;
defparam \macro_inst|controller|sm_pwm|pwmCnt[4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmCnt[4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[4] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmCnt[5] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|Add0~9 ),
	.Qin(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|pwmUpdateTrigger~q_X59_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Add0~10_combout ),
	.Cout(\macro_inst|controller|sm_pwm|Add0~11 ),
	.Q(\macro_inst|controller|sm_pwm|pwmCnt [5]));
defparam \macro_inst|controller|sm_pwm|pwmCnt[5] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmCnt[5] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmCnt[5] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmCnt[5] .mask = 16'h3C3F;
defparam \macro_inst|controller|sm_pwm|pwmCnt[5] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmCnt[5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[5] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmCnt[6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|Add0~11 ),
	.Qin(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|pwmUpdateTrigger~q_X59_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|Add0~12_combout ),
	.Cout(\macro_inst|controller|sm_pwm|Add0~13 ),
	.Q(\macro_inst|controller|sm_pwm|pwmCnt [6]));
defparam \macro_inst|controller|sm_pwm|pwmCnt[6] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmCnt[6] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmCnt[6] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmCnt[6] .mask = 16'hC30C;
defparam \macro_inst|controller|sm_pwm|pwmCnt[6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmCnt[6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[6] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[6] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmCnt[7] (
	.A(\macro_inst|controller|sm_pwm|Add0~14_combout ),
	.B(vcc),
	.C(\macro_inst|controller|sm_pwm|Equal1~1_combout ),
	.D(\macro_inst|controller|sm_pwm|Equal1~0_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|pwmUpdateTrigger~q_X59_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmCnt~0_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmCnt [7]));
defparam \macro_inst|controller|sm_pwm|pwmCnt[7] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmCnt[7] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmCnt[7] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmCnt[7] .mask = 16'h0AAA;
defparam \macro_inst|controller|sm_pwm|pwmCnt[7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmCnt[7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X59_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[0][0]~49_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][0] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[0][0] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[0][0] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[0][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[0][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan1~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(SyncReset_X59_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan1~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][10] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[0][10] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[0][10] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[0][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[0][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[0][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan1~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(SyncReset_X59_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan1~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][11] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[0][11] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[0][11] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[0][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[0][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[0][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan1~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(SyncReset_X59_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan1~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][12] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[0][12] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[0][12] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[0][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[0][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][13] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[0][13]~q ),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan1~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(SyncReset_X59_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan1~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][13] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[0][13] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[0][13] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[0][13] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[0][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[0][14]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan1~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(SyncReset_X59_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y9_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan1~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][14] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[0][14] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[0][14] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[0][14] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[0][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][15] (
	.A(\macro_inst|controller|sm_pwm|LessThan2~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[0][7]~q ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X61_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ),
	.SyncReset(SyncReset_X61_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y11_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~216_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][15] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[0][15] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[0][15] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[0][15] .mask = 16'h77F0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[0][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan2~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X61_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ),
	.SyncReset(SyncReset_X61_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan2~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][1] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[0][1] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[0][1] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[0][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[0][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[0][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan2~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X61_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ),
	.SyncReset(SyncReset_X61_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan2~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][2] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[0][2] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[0][2] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[0][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[0][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[0][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan2~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X61_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ),
	.SyncReset(SyncReset_X61_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan2~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][3] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[0][3] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[0][3] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[0][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[0][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[0][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan2~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X61_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ),
	.SyncReset(SyncReset_X61_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan2~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][4] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[0][4] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[0][4] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[0][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[0][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X60_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[0][5]~48_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][5] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[0][5] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[0][5] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[0][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[0][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan2~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X61_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y11_SIG ),
	.SyncReset(SyncReset_X61_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y11_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan2~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][6] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[0][6] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[0][6] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[0][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[0][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][7] (
	.A(\macro_inst|controller|sm_pwm|pwmList[31][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(SyncReset_X59_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan64~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][7] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[0][7] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[0][7] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[0][7] .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|pwmList[0][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][7] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[0][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(SyncReset_X59_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan1~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][8] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[0][8] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[0][8] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[0][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[0][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[0][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[0][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan1~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[0][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~49_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(SyncReset_X59_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan1~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[0][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[0][9] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[0][9] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[0][9] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[0][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[0][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[0][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[0][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][0] (
	.A(vcc),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[0] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X62_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[10][0]~87_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][0] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[10][0] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[10][0] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[10][0] .mask = 16'h0F0F;
defparam \macro_inst|controller|sm_pwm|pwmList[10][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[10][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan21~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X61_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y10_SIG ),
	.SyncReset(SyncReset_X61_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan21~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][10] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[10][10] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[10][10] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[10][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[10][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][11] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[10][11]~q ),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan21~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X61_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y10_SIG ),
	.SyncReset(SyncReset_X61_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan21~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][11] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[10][11] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[10][11] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[10][11] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[10][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[10][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan21~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X61_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y10_SIG ),
	.SyncReset(SyncReset_X61_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan21~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][12] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[10][12] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[10][12] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[10][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[10][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[10][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X62_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(SyncReset_X62_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan22~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][13] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[10][13] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[10][13] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[10][13] .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|pwmList[10][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][14] (
	.A(\macro_inst|controller|sm_pwm|pwmList[10][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan22~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X62_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(SyncReset_X62_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan22~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][14] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[10][14] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[10][14] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[10][14] .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|pwmList[10][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][14] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][15] (
	.A(\macro_inst|controller|sm_pwm|LessThan22~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[10][7]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X62_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(SyncReset_X62_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y10_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~254_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][15] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[10][15] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[10][15] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[10][15] .mask = 16'h74FC;
defparam \macro_inst|controller|sm_pwm|pwmList[10][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[10][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan22~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X62_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(SyncReset_X62_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan22~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][1] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[10][1] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[10][1] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[10][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[10][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[10][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan22~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X62_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(SyncReset_X62_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan22~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][2] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[10][2] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[10][2] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[10][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[10][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[10][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan22~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X62_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(SyncReset_X62_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan22~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][3] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[10][3] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[10][3] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[10][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[10][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[10][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan22~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X62_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(SyncReset_X62_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan22~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][4] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[10][4] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[10][4] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[10][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[10][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X62_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[10][5]~86_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][5] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[10][5] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[10][5] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[10][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[10][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[10][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan22~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X62_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(SyncReset_X62_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y10_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan22~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][6] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[10][6] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[10][6] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[10][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[10][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][7] (
	.A(\macro_inst|controller|sm_pwm|pwmList[10][15]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|LessThan21~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X62_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y10_SIG ),
	.SyncReset(SyncReset_X62_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y10_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~206_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][7] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[10][7] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[10][7] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[10][7] .mask = 16'h8BCF;
defparam \macro_inst|controller|sm_pwm|pwmList[10][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][8] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[8] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X61_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[10][8]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][8] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[10][8] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[10][8] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[10][8] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[10][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][8] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][8] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[10][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[10][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan21~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[10][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~74_combout_X61_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y10_SIG ),
	.SyncReset(SyncReset_X61_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan21~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[10][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[10][9] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[10][9] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[10][9] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[10][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[10][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[10][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[10][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X62_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[11][0]~39_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][0] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[11][0] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[11][0] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[11][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[11][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan23~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan23~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][10] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[11][10] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[11][10] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[11][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[11][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[11][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan23~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan23~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][11] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[11][11] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[11][11] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[11][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[11][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][12] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[11][12]~q ),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan23~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan23~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][12] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[11][12] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[11][12] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[11][12] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[11][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][13] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[11][13]~q ),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan23~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan23~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][13] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[11][13] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[11][13] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[11][13] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[11][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[11][14]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan23~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan23~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][14] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[11][14] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[11][14] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[11][14] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[11][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][15] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[11][7]~q ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|LessThan24~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X61_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(SyncReset_X61_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~110_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][15] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[11][15] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[11][15] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[11][15] .mask = 16'h72FA;
defparam \macro_inst|controller|sm_pwm|pwmList[11][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][1] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [8]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[8]~8_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][1] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[11][1] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[11][1] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][1] .mask = 16'hCC00;
defparam \macro_inst|controller|sm_pwm|pwmList[11][1] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][1] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[11][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan24~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X62_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ),
	.SyncReset(SyncReset_X62_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan24~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][2] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[11][2] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[11][2] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[11][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[11][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[11][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan24~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X62_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ),
	.SyncReset(SyncReset_X62_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan24~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][3] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[11][3] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[11][3] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[11][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[11][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[11][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan24~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X62_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ),
	.SyncReset(SyncReset_X62_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan24~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][4] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[11][4] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[11][4] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[11][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[11][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][5] (
	.A(vcc),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[5] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X62_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[11][5]~38_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][5] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[11][5] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[11][5] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[11][5] .mask = 16'h0F0F;
defparam \macro_inst|controller|sm_pwm|pwmList[11][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[11][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan24~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X62_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y2_SIG ),
	.SyncReset(SyncReset_X62_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y2_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan24~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][6] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[11][6] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[11][6] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[11][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[11][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][7] (
	.A(\macro_inst|controller|sm_pwm|pwmList[11][15]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan23~12_combout ),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X61_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y4_SIG ),
	.SyncReset(SyncReset_X61_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~62_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][7] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[11][7] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[11][7] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[11][7] .mask = 16'hBB0F;
defparam \macro_inst|controller|sm_pwm|pwmList[11][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][8] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[11][8]~q ),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan23~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][8] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[11][8] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[11][8] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[11][8] .mask = 16'h0044;
defparam \macro_inst|controller|sm_pwm|pwmList[11][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[11][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[11][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan23~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[11][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~44_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan23~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[11][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[11][9] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[11][9] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[11][9] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[11][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[11][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[11][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[11][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X58_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[12][0]~89_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][0] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[12][0] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[12][0] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[12][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[12][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[12][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan25~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X57_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ),
	.SyncReset(SyncReset_X57_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan25~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][10] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[12][10] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[12][10] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[12][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[12][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[12][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan25~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X57_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ),
	.SyncReset(SyncReset_X57_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan25~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][11] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[12][11] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[12][11] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[12][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[12][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[12][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan26~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X58_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(SyncReset_X58_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan26~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][12] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[12][12] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[12][12] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[12][12] .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|pwmList[12][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[12][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan25~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X57_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ),
	.SyncReset(SyncReset_X57_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan25~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][13] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[12][13] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[12][13] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[12][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[12][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[12][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan25~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X57_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ),
	.SyncReset(SyncReset_X57_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y11_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan25~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][14] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[12][14] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[12][14] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[12][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[12][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][15] (
	.A(\macro_inst|controller|sm_pwm|LessThan26~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[12][7]~q ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X58_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(SyncReset_X58_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y11_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~256_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][15] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[12][15] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[12][15] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[12][15] .mask = 16'h77F0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[12][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan26~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X58_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(SyncReset_X58_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan26~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][1] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[12][1] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[12][1] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[12][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[12][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[12][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan26~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X58_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(SyncReset_X58_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan26~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][2] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[12][2] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[12][2] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[12][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[12][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[12][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan26~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X58_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(SyncReset_X58_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan26~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][3] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[12][3] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[12][3] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[12][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[12][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[12][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan26~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X58_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(SyncReset_X58_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan26~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][4] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[12][4] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[12][4] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[12][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[12][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][5] (
	.A(vcc),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[5] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X58_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[12][5]~88_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][5] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[12][5] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[12][5] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][5] .mask = 16'h0F0F;
defparam \macro_inst|controller|sm_pwm|pwmList[12][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[12][6]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan26~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X58_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(SyncReset_X58_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y11_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan26~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][6] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[12][6] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[12][6] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[12][6] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[12][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][7] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[12][15]~q ),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|LessThan25~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X58_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(SyncReset_X58_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y11_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~208_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][7] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[12][7] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[12][7] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[12][7] .mask = 16'h8DAF;
defparam \macro_inst|controller|sm_pwm|pwmList[12][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[12][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X57_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ),
	.SyncReset(SyncReset_X57_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan25~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][8] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[12][8] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[12][8] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[12][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[12][9] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[12][0]~q ),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[12][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~76_combout_X58_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y11_SIG ),
	.SyncReset(SyncReset_X58_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan26~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[12][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[12][9] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[12][9] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[12][9] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[12][9] .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|pwmList[12][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[12][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[12][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[13][0]~41_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][0] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[13][0] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[13][0] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[13][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[13][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan27~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(SyncReset_X59_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan27~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][10] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[13][10] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[13][10] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[13][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[13][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][11] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[13][11]~q ),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan27~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(SyncReset_X59_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan27~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][11] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[13][11] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[13][11] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[13][11] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[13][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][12] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[13][12]~q ),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan27~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(SyncReset_X59_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan27~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][12] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[13][12] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[13][12] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[13][12] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[13][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[13][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan27~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(SyncReset_X59_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan27~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][13] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[13][13] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[13][13] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[13][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[13][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[13][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan27~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(SyncReset_X59_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y8_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan27~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][14] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[13][14] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[13][14] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[13][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[13][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][15] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [10]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y4_SIG ),
	.SyncReset(SyncReset_X59_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y4_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[10]~10_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][15] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[13][15] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[13][15] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[13][15] .mask = 16'hCC00;
defparam \macro_inst|controller|sm_pwm|pwmList[13][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[13][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan28~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X58_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y4_SIG ),
	.SyncReset(SyncReset_X58_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan28~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][1] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[13][1] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[13][1] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[13][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[13][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][2] (
	.A(\macro_inst|ahb_add_reg [1]),
	.B(\macro_inst|ahb_add_reg [5]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(\macro_inst|ahb_add_reg [6]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y4_SIG ),
	.SyncReset(SyncReset_X59_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~10_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][2] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[13][2] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[13][2] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[13][2] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[13][2] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][2] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[13][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan28~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X58_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y4_SIG ),
	.SyncReset(SyncReset_X58_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan28~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][3] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[13][3] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[13][3] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[13][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[13][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[13][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan28~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X58_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y4_SIG ),
	.SyncReset(SyncReset_X58_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan28~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][4] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[13][4] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[13][4] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[13][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[13][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[13][5]~40_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][5] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[13][5] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[13][5] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[13][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[13][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[13][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan28~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X58_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y4_SIG ),
	.SyncReset(SyncReset_X58_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan28~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][6] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[13][6] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[13][6] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[13][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[13][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][7] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [14]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y4_SIG ),
	.SyncReset(SyncReset_X59_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y4_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[14]~14_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][7] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[13][7] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[13][7] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[13][7] .mask = 16'hCC00;
defparam \macro_inst|controller|sm_pwm|pwmList[13][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[13][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(SyncReset_X59_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan27~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][8] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[13][8] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[13][8] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[13][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[13][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[13][9] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[13][9]~q ),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan27~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[13][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~45_combout_X59_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y8_SIG ),
	.SyncReset(SyncReset_X59_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan27~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[13][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[13][9] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[13][9] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[13][9] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[13][9] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[13][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[13][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[13][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][0] (
	.A(vcc),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[0] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X62_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[14][0]~91_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][0] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[14][0] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[14][0] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[14][0] .mask = 16'h0F0F;
defparam \macro_inst|controller|sm_pwm|pwmList[14][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[14][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan29~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X61_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ),
	.SyncReset(SyncReset_X61_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan29~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][10] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[14][10] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[14][10] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[14][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[14][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[14][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan29~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X61_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ),
	.SyncReset(SyncReset_X61_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan29~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][11] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[14][11] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[14][11] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[14][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[14][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][12] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[14][12]~q ),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan29~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X61_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ),
	.SyncReset(SyncReset_X61_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan29~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][12] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[14][12] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[14][12] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[14][12] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[14][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][13] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[14][13]~q ),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan29~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X61_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ),
	.SyncReset(SyncReset_X61_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan29~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][13] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[14][13] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[14][13] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[14][13] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[14][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[14][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan29~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X61_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ),
	.SyncReset(SyncReset_X61_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan29~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][14] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[14][14] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[14][14] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[14][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[14][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[14][7]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan30~12_combout ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X62_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ),
	.SyncReset(SyncReset_X62_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~258_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][15] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[14][15] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[14][15] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[14][15] .mask = 16'h77F0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][1] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[14][1]~q ),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan30~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X62_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ),
	.SyncReset(SyncReset_X62_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan30~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][1] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[14][1] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[14][1] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[14][1] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[14][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[14][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan30~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X62_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ),
	.SyncReset(SyncReset_X62_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan30~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][2] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[14][2] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[14][2] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[14][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[14][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[14][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan30~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X62_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ),
	.SyncReset(SyncReset_X62_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan30~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][3] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[14][3] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[14][3] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[14][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[14][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[14][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan30~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X62_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ),
	.SyncReset(SyncReset_X62_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan30~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][4] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[14][4] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[14][4] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[14][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[14][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X62_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[14][5]~90_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][5] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[14][5] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[14][5] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[14][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[14][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[14][6]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan30~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X62_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ),
	.SyncReset(SyncReset_X62_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan30~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][6] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[14][6] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[14][6] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[14][6] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[14][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][7] (
	.A(\macro_inst|controller|sm_pwm|pwmList[14][15]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan29~12_combout ),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X62_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y3_SIG ),
	.SyncReset(SyncReset_X62_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~210_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][7] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[14][7] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[14][7] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[14][7] .mask = 16'hBB0F;
defparam \macro_inst|controller|sm_pwm|pwmList[14][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[14][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X61_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ),
	.SyncReset(SyncReset_X61_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan29~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][8] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[14][8] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[14][8] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[14][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[14][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[14][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan29~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[14][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~77_combout_X61_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ),
	.SyncReset(SyncReset_X61_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan29~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[14][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[14][9] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[14][9] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[14][9] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[14][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[14][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[14][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[14][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][0] (
	.A(vcc),
	.B(\rv32.mem_ahb_hwdata[0] ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X60_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[15][0]~43_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][0] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[15][0] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[15][0] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[15][0] .mask = 16'h3333;
defparam \macro_inst|controller|sm_pwm|pwmList[15][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[15][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan31~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X61_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ),
	.SyncReset(SyncReset_X61_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan31~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][10] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[15][10] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[15][10] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[15][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[15][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[15][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan31~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X61_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ),
	.SyncReset(SyncReset_X61_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan31~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][11] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[15][11] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[15][11] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[15][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[15][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][12] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[15][12]~q ),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan31~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X61_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ),
	.SyncReset(SyncReset_X61_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan31~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][12] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[15][12] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[15][12] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[15][12] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[15][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][13] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[15][13]~q ),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan31~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X61_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ),
	.SyncReset(SyncReset_X61_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan31~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][13] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[15][13] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[15][13] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[15][13] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[15][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][14] (
	.A(\macro_inst|controller|sm_pwm|pwmList[15][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan32~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X60_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y7_SIG ),
	.SyncReset(SyncReset_X60_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan32~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][14] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[15][14] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[15][14] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[15][14] .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|pwmList[15][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][14] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[15][7]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan32~12_combout ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X61_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ),
	.SyncReset(SyncReset_X61_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~114_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][15] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[15][15] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[15][15] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][15] .mask = 16'h77F0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[15][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan32~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X60_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y7_SIG ),
	.SyncReset(SyncReset_X60_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan32~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][1] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[15][1] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[15][1] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[15][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[15][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[15][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan32~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X60_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y7_SIG ),
	.SyncReset(SyncReset_X60_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan32~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][2] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[15][2] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[15][2] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[15][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[15][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[15][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan32~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X60_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y7_SIG ),
	.SyncReset(SyncReset_X60_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan32~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][3] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[15][3] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[15][3] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[15][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[15][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[15][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan32~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X60_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y7_SIG ),
	.SyncReset(SyncReset_X60_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan32~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][4] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[15][4] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[15][4] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[15][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[15][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X60_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[15][5]~42_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][5] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[15][5] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[15][5] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[15][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[15][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan32~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X60_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y7_SIG ),
	.SyncReset(SyncReset_X60_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan32~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][6] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[15][6] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[15][6] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[15][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[15][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][7] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[15][0]~q ),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X60_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y7_SIG ),
	.SyncReset(SyncReset_X60_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan32~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][7] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[15][7] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[15][7] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[15][7] .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|pwmList[15][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][7] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[15][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X61_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ),
	.SyncReset(SyncReset_X61_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan31~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][8] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[15][8] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[15][8] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[15][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[15][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[15][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[15][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan31~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[15][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~46_combout_X61_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y7_SIG ),
	.SyncReset(SyncReset_X61_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan31~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[15][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[15][9] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[15][9] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[15][9] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[15][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[15][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[15][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[15][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X59_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[16][0]~93_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][0] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[16][0] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[16][0] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[16][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[16][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[16][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan33~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X56_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y2_SIG ),
	.SyncReset(SyncReset_X56_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan33~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][10] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[16][10] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[16][10] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[16][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[16][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][11] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[16][11]~q ),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan33~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X56_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y2_SIG ),
	.SyncReset(SyncReset_X56_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan33~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][11] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[16][11] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[16][11] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[16][11] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[16][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[16][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan33~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X56_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y2_SIG ),
	.SyncReset(SyncReset_X56_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan33~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][12] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[16][12] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[16][12] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[16][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[16][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][13] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[16][13]~q ),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan33~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X56_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y2_SIG ),
	.SyncReset(SyncReset_X56_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan33~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][13] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[16][13] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[16][13] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[16][13] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[16][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][14] (
	.A(\macro_inst|controller|sm_pwm|pwmList[16][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan34~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X59_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ),
	.SyncReset(SyncReset_X59_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan34~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][14] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[16][14] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[16][14] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[16][14] .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|pwmList[16][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][14] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][15] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[16][7]~q ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|LessThan34~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X59_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ),
	.SyncReset(SyncReset_X59_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y2_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~260_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][15] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[16][15] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[16][15] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[16][15] .mask = 16'h72FA;
defparam \macro_inst|controller|sm_pwm|pwmList[16][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[16][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan34~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X59_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ),
	.SyncReset(SyncReset_X59_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan34~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][1] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[16][1] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[16][1] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[16][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][2] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.B(\macro_inst|controller|sm_pwm|pwmList[16][2]~q ),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan34~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X59_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ),
	.SyncReset(SyncReset_X59_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan34~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][2] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[16][2] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[16][2] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[16][2] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[16][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[16][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan34~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X59_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ),
	.SyncReset(SyncReset_X59_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan34~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][3] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[16][3] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[16][3] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[16][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[16][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[16][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan34~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X59_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ),
	.SyncReset(SyncReset_X59_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan34~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][4] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[16][4] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[16][4] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[16][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[16][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X59_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[16][5]~92_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][5] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[16][5] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[16][5] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[16][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[16][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[16][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan34~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X59_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ),
	.SyncReset(SyncReset_X59_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y2_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan34~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][6] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[16][6] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[16][6] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[16][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[16][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][7] (
	.A(\macro_inst|controller|sm_pwm|LessThan33~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[16][15]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X59_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y2_SIG ),
	.SyncReset(SyncReset_X59_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y2_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~212_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][7] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[16][7] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[16][7] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[16][7] .mask = 16'hCF47;
defparam \macro_inst|controller|sm_pwm|pwmList[16][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[16][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X56_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y2_SIG ),
	.SyncReset(SyncReset_X56_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan33~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][8] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[16][8] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[16][8] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[16][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[16][9] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[16][9]~q ),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan33~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[16][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~78_combout_X56_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y2_SIG ),
	.SyncReset(SyncReset_X56_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan33~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[16][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[16][9] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[16][9] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[16][9] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][9] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[16][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[16][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[16][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[17][0]~45_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][0] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[17][0] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][0] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[17][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[17][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[17][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan35~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(SyncReset_X61_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan35~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][10] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[17][10] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][10] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[17][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[17][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[17][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan35~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(SyncReset_X61_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan35~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][11] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[17][11] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][11] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[17][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[17][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[17][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan35~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(SyncReset_X61_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan35~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][12] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[17][12] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][12] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[17][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[17][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[17][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan35~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(SyncReset_X61_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan35~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][13] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[17][13] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][13] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[17][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[17][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[17][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan35~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(SyncReset_X61_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan35~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][14] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[17][14] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][14] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[17][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[17][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][15] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[15] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X62_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[17][15]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][15] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[17][15] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][15] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[17][15] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[17][15] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][15] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[17][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan36~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X62_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y1_SIG ),
	.SyncReset(SyncReset_X62_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan36~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][1] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[17][1] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][1] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[17][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[17][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][2] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.B(\macro_inst|controller|sm_pwm|pwmList[17][2]~q ),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan36~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X62_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y1_SIG ),
	.SyncReset(SyncReset_X62_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan36~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][2] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[17][2] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][2] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[17][2] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[17][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[17][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan36~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X62_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y1_SIG ),
	.SyncReset(SyncReset_X62_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan36~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][3] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[17][3] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][3] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[17][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[17][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[17][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan36~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X62_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y1_SIG ),
	.SyncReset(SyncReset_X62_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan36~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][4] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[17][4] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][4] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[17][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[17][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][5] (
	.A(vcc),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[5] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[17][5]~44_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][5] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[17][5] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][5] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][5] .mask = 16'h0F0F;
defparam \macro_inst|controller|sm_pwm|pwmList[17][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][6] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[17][6]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan36~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X62_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y1_SIG ),
	.SyncReset(SyncReset_X62_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y1_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan36~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][6] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[17][6] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][6] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[17][6] .mask = 16'h5F05;
defparam \macro_inst|controller|sm_pwm|pwmList[17][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X62_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[17][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][7] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[17][7] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][7] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[17][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[17][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[17][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(SyncReset_X61_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan35~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][8] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[17][8] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][8] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[17][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[17][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[17][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[17][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan35~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[17][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~81_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(SyncReset_X61_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan35~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[17][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[17][9] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[17][9] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][9] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[17][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[17][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[17][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[17][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X54_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[18][0]~95_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][0] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[18][0] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[18][0] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[18][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[18][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[18][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan37~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan37~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][10] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[18][10] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[18][10] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[18][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[18][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[18][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan37~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan37~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][11] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[18][11] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[18][11] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[18][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[18][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][12] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[18][12]~q ),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan37~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan37~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][12] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[18][12] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[18][12] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[18][12] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[18][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][13] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[18][13]~q ),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan37~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan37~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][13] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[18][13] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[18][13] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[18][13] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[18][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[18][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan37~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan37~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][14] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[18][14] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[18][14] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[18][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[18][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][15] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|LessThan38~12_combout ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[18][7]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X54_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ),
	.SyncReset(SyncReset_X54_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~262_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][15] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[18][15] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[18][15] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[18][15] .mask = 16'h72FA;
defparam \macro_inst|controller|sm_pwm|pwmList[18][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][1] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[18][1]~q ),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan38~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X54_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ),
	.SyncReset(SyncReset_X54_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan38~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][1] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[18][1] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[18][1] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][1] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[18][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[18][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan38~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X54_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ),
	.SyncReset(SyncReset_X54_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan38~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][2] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[18][2] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[18][2] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[18][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[18][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[18][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan38~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X54_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ),
	.SyncReset(SyncReset_X54_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan38~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][3] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[18][3] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[18][3] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[18][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[18][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[18][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan38~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X54_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ),
	.SyncReset(SyncReset_X54_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan38~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][4] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[18][4] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[18][4] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[18][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[18][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X54_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[18][5]~94_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][5] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[18][5] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[18][5] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[18][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[18][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[18][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan38~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X54_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ),
	.SyncReset(SyncReset_X54_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan38~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][6] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[18][6] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[18][6] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[18][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[18][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X54_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[18][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][7] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[18][7] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[18][7] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[18][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[18][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][8] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [1]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[1]~1_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][8] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[18][8] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[18][8] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[18][8] .mask = 16'hCC00;
defparam \macro_inst|controller|sm_pwm|pwmList[18][8] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][8] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[18][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[18][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan37~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[18][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~79_combout_X58_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y6_SIG ),
	.SyncReset(SyncReset_X58_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan37~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[18][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[18][9] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[18][9] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[18][9] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[18][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[18][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[18][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[18][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X62_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[19][0]~47_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][0] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[19][0] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[19][0] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[19][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[19][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[19][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan39~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan39~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][10] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[19][10] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[19][10] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[19][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[19][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[19][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan39~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan39~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][11] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[19][11] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[19][11] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[19][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[19][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[19][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan39~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan39~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][12] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[19][12] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[19][12] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[19][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[19][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][13] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[19][13]~q ),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan39~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan39~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][13] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[19][13] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[19][13] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[19][13] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[19][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[19][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan39~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan39~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][14] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[19][14] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[19][14] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[19][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[19][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][15] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[15] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X62_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[19][15]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][15] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[19][15] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[19][15] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[19][15] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[19][15] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][15] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[19][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan40~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X62_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y4_SIG ),
	.SyncReset(SyncReset_X62_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan40~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][1] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[19][1] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[19][1] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[19][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[19][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[19][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan40~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X62_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y4_SIG ),
	.SyncReset(SyncReset_X62_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan40~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][2] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[19][2] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[19][2] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[19][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[19][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[19][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan40~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X62_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y4_SIG ),
	.SyncReset(SyncReset_X62_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan40~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][3] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[19][3] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[19][3] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[19][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[19][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[19][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan40~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X62_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y4_SIG ),
	.SyncReset(SyncReset_X62_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan40~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][4] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[19][4] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[19][4] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[19][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[19][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][5] (
	.A(vcc),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[5] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X62_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[19][5]~46_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][5] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[19][5] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[19][5] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][5] .mask = 16'h0F0F;
defparam \macro_inst|controller|sm_pwm|pwmList[19][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[19][6]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan40~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X62_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y4_SIG ),
	.SyncReset(SyncReset_X62_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan40~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][6] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[19][6] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[19][6] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[19][6] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[19][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X62_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[19][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][7] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[19][7] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[19][7] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[19][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[19][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[19][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan39~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][8] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[19][8] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[19][8] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[19][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[19][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[19][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[19][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan39~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[19][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~47_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan39~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[19][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[19][9] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[19][9] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[19][9] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[19][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[19][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[19][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[19][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X59_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[1][0]~1_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][0] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[1][0] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[1][0] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[1][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[1][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[1][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan3~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan3~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][10] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[1][10] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[1][10] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[1][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[1][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[1][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan3~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan3~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][11] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[1][11] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[1][11] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[1][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[1][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[1][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan3~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan3~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][12] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[1][12] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[1][12] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[1][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[1][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[1][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan3~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan3~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][13] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[1][13] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[1][13] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[1][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[1][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[1][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan3~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan3~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][14] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[1][14] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[1][14] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[1][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[1][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][15] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[1][7]~q ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|LessThan4~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~72_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][15] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[1][15] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[1][15] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[1][15] .mask = 16'h72FA;
defparam \macro_inst|controller|sm_pwm|pwmList[1][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[1][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan4~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X59_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ),
	.SyncReset(SyncReset_X59_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan4~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][1] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[1][1] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[1][1] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[1][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[1][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[1][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan4~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X59_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ),
	.SyncReset(SyncReset_X59_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan4~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][2] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[1][2] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[1][2] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[1][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[1][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][3] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[1][3]~q ),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan4~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X59_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ),
	.SyncReset(SyncReset_X59_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan4~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][3] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[1][3] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[1][3] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[1][3] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[1][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[1][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan4~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X59_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ),
	.SyncReset(SyncReset_X59_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan4~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][4] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[1][4] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[1][4] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[1][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[1][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X59_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[1][5]~0_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][5] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[1][5] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[1][5] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[1][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[1][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[1][6]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan4~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X59_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ),
	.SyncReset(SyncReset_X59_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan4~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][6] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[1][6] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[1][6] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[1][6] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[1][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][7] (
	.A(\macro_inst|controller|sm_pwm|pwmList[1][15]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|LessThan3~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~24_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][7] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[1][7] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[1][7] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[1][7] .mask = 16'h8BCF;
defparam \macro_inst|controller|sm_pwm|pwmList[1][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[1][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan3~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][8] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[1][8] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[1][8] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[1][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[1][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[1][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[1][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan3~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[1][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~11_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan3~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[1][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[1][9] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[1][9] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[1][9] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[1][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[1][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[1][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[1][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[20][0]~53_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][0] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[20][0] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[20][0] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[20][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[20][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[20][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan41~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(SyncReset_X60_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan41~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][10] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[20][10] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[20][10] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[20][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[20][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][11] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[20][11]~q ),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan41~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(SyncReset_X60_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan41~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][11] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[20][11] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[20][11] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[20][11] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[20][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[20][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan41~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(SyncReset_X60_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan41~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][12] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[20][12] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[20][12] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[20][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[20][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[20][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan41~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(SyncReset_X60_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan41~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][13] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[20][13] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[20][13] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[20][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[20][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[20][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan41~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(SyncReset_X60_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y2_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan41~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][14] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[20][14] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[20][14] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[20][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[20][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][15] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[15] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X54_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[20][15]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][15] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[20][15] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[20][15] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[20][15] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[20][15] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][15] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[20][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan42~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X54_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y2_SIG ),
	.SyncReset(SyncReset_X54_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan42~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][1] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[20][1] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[20][1] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[20][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[20][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[20][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan42~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X54_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y2_SIG ),
	.SyncReset(SyncReset_X54_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan42~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][2] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[20][2] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[20][2] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[20][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[20][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[20][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan42~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X54_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y2_SIG ),
	.SyncReset(SyncReset_X54_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan42~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][3] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[20][3] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[20][3] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[20][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[20][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[20][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan42~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X54_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y2_SIG ),
	.SyncReset(SyncReset_X54_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan42~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][4] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[20][4] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[20][4] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[20][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[20][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X54_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[20][5]~52_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][5] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[20][5] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[20][5] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[20][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[20][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][6] (
	.A(\macro_inst|controller|sm_pwm|pwmList[20][6]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan42~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X54_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y2_SIG ),
	.SyncReset(SyncReset_X54_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X54_Y2_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan42~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][6] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[20][6] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[20][6] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[20][6] .mask = 16'h2B2B;
defparam \macro_inst|controller|sm_pwm|pwmList[20][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X54_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[20][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][7] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[20][7] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[20][7] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[20][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[20][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[20][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(SyncReset_X60_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan41~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][8] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[20][8] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[20][8] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[20][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[20][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[20][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan41~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[20][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~52_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(SyncReset_X60_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan41~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[20][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[20][9] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[20][9] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[20][9] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[20][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[20][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[20][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[20][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X57_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[21][0]~5_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][0] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[21][0] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[21][0] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[21][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[21][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][10] (
	.A(\macro_inst|ahb_add_reg [1]),
	.B(\macro_inst|ahb_add_reg [5]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(\macro_inst|ahb_add_reg [6]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X57_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ),
	.SyncReset(SyncReset_X57_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y2_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~16_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][10] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[21][10] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[21][10] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[21][10] .mask = 16'h0088;
defparam \macro_inst|controller|sm_pwm|pwmList[21][10] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][10] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][11] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[21][11]~q ),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan43~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X56_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y2_SIG ),
	.SyncReset(SyncReset_X56_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan43~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][11] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[21][11] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[21][11] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[21][11] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[21][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[21][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan44~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X57_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ),
	.SyncReset(SyncReset_X57_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan44~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][12] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[21][12] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[21][12] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[21][12] .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|pwmList[21][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][13] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[21][13]~q ),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan43~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X56_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y2_SIG ),
	.SyncReset(SyncReset_X56_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan43~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][13] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[21][13] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[21][13] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[21][13] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[21][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][14] (
	.A(\macro_inst|controller|sm_pwm|pwmList[21][14]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan43~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X56_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y2_SIG ),
	.SyncReset(SyncReset_X56_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y2_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan43~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][14] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[21][14] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[21][14] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[21][14] .mask = 16'h2B2B;
defparam \macro_inst|controller|sm_pwm|pwmList[21][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[21][7]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan44~12_combout ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X57_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ),
	.SyncReset(SyncReset_X57_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y2_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~76_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][15] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[21][15] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[21][15] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][15] .mask = 16'h77F0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[21][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan44~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X57_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ),
	.SyncReset(SyncReset_X57_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan44~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][1] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[21][1] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[21][1] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[21][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[21][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[21][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan44~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X57_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ),
	.SyncReset(SyncReset_X57_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan44~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][2] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[21][2] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[21][2] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[21][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[21][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[21][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan44~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X57_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ),
	.SyncReset(SyncReset_X57_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan44~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][3] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[21][3] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[21][3] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[21][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[21][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[21][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan44~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X57_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ),
	.SyncReset(SyncReset_X57_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan44~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][4] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[21][4] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[21][4] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[21][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[21][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X56_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[21][5]~4_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][5] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[21][5] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[21][5] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[21][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[21][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[21][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan44~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X57_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ),
	.SyncReset(SyncReset_X57_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y2_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan44~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][6] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[21][6] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[21][6] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[21][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[21][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][7] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[21][0]~q ),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X57_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y2_SIG ),
	.SyncReset(SyncReset_X57_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan44~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][7] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[21][7] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[21][7] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[21][7] .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|pwmList[21][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][7] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[21][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X56_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y2_SIG ),
	.SyncReset(SyncReset_X56_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan43~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][8] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[21][8] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[21][8] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[21][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[21][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[21][9] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[21][9]~q ),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan43~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[21][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~17_combout_X56_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y2_SIG ),
	.SyncReset(SyncReset_X56_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan43~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[21][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[21][9] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[21][9] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[21][9] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[21][9] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[21][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[21][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[21][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X56_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[22][0]~55_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][0] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][0] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[22][0] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[22][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[22][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[22][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan45~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(SyncReset_X58_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan45~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][10] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][10] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][10] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[22][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[22][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan45~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(SyncReset_X58_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan45~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][11] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][11] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][11] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[22][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[22][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[22][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan45~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(SyncReset_X58_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan45~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][12] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][12] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][12] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[22][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[22][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[22][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan45~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(SyncReset_X58_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan45~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][13] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][13] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][13] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[22][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[22][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[22][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan45~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(SyncReset_X58_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y1_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan45~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][14] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][14] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][14] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[22][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[22][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[22][7]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|LessThan46~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X56_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ),
	.SyncReset(SyncReset_X56_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y1_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~222_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][15] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][15] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[22][15] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[22][15] .mask = 16'h74FC;
defparam \macro_inst|controller|sm_pwm|pwmList[22][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][1] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[22][1]~q ),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan46~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X56_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ),
	.SyncReset(SyncReset_X56_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan46~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][1] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][1] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[22][1] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][1] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[22][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[22][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan46~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X56_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ),
	.SyncReset(SyncReset_X56_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan46~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][2] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][2] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[22][2] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[22][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[22][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[22][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan46~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X56_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ),
	.SyncReset(SyncReset_X56_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan46~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][3] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][3] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[22][3] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[22][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[22][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[22][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan46~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X56_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ),
	.SyncReset(SyncReset_X56_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan46~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][4] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][4] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[22][4] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[22][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[22][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X56_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[22][5]~54_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][5] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][5] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[22][5] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[22][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[22][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[22][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan46~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X56_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ),
	.SyncReset(SyncReset_X56_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y1_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan46~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][6] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][6] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[22][6] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[22][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[22][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][7] (
	.A(\macro_inst|controller|sm_pwm|pwmList[22][15]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|LessThan45~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X56_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y1_SIG ),
	.SyncReset(SyncReset_X56_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y1_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~174_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][7] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][7] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[22][7] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][7] .mask = 16'h8BCF;
defparam \macro_inst|controller|sm_pwm|pwmList[22][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[22][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(SyncReset_X58_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan45~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][8] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][8] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][8] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[22][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[22][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[22][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[22][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan45~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[22][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~54_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(SyncReset_X58_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan45~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[22][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[22][9] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[22][9] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][9] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[22][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[22][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[22][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[22][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X62_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[23][0]~7_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][0] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[23][0] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[23][0] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[23][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][10] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[23][14]~q ),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan47~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan47~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][10] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[23][10] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[23][10] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[23][10] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[23][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][10] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[23][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan47~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan47~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][11] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[23][11] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[23][11] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[23][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[23][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[23][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan47~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan47~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][12] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[23][12] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[23][12] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[23][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[23][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[23][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan47~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][13] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[23][13] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[23][13] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[23][13] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[23][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][14] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[23][11]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan47~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan47~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][14] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[23][14] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[23][14] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[23][14] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[23][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][14] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][15] (
	.A(\macro_inst|controller|sm_pwm|LessThan47~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[23][7]~q ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~30_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][15] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[23][15] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[23][15] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[23][15] .mask = 16'hF533;
defparam \macro_inst|controller|sm_pwm|pwmList[23][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[23][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan48~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X62_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y6_SIG ),
	.SyncReset(SyncReset_X62_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan48~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][1] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[23][1] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[23][1] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[23][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[23][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[23][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan48~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X62_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y6_SIG ),
	.SyncReset(SyncReset_X62_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan48~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][2] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[23][2] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[23][2] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[23][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[23][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][3] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[23][3]~q ),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan48~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X62_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y6_SIG ),
	.SyncReset(SyncReset_X62_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan48~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][3] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[23][3] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[23][3] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[23][3] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[23][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[23][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan48~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X62_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y6_SIG ),
	.SyncReset(SyncReset_X62_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan48~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][4] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[23][4] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[23][4] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[23][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[23][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][5] (
	.A(vcc),
	.B(\rv32.mem_ahb_hwdata[5] ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X62_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[23][5]~6_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][5] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[23][5] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[23][5] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[23][5] .mask = 16'h3333;
defparam \macro_inst|controller|sm_pwm|pwmList[23][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][6] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[23][6]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan48~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X62_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y6_SIG ),
	.SyncReset(SyncReset_X62_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y6_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan48~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][6] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[23][6] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[23][6] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[23][6] .mask = 16'h5F05;
defparam \macro_inst|controller|sm_pwm|pwmList[23][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X62_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[23][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][7] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[23][7] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[23][7] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[23][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[23][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[23][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan47~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan47~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][8] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[23][8] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[23][8] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[23][8] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[23][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[23][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[23][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan47~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[23][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~20_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan47~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[23][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[23][9] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[23][9] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[23][9] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[23][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[23][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[23][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[23][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X56_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[24][0]~57_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][0] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[24][0] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][0] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[24][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[24][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[24][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan49~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(SyncReset_X58_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan49~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][10] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[24][10] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][10] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[24][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[24][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[24][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan49~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(SyncReset_X58_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan49~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][11] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[24][11] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][11] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[24][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[24][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][12] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[24][12]~q ),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan49~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(SyncReset_X58_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan49~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][12] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[24][12] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][12] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[24][12] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[24][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[24][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan49~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(SyncReset_X58_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan49~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][13] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[24][13] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][13] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[24][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[24][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[24][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan49~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(SyncReset_X58_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y9_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan49~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][14] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[24][14] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][14] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[24][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[24][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[24][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan50~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X56_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y9_SIG ),
	.SyncReset(SyncReset_X56_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan50~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][15] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[24][15] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][15] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[24][15] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[24][15] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][15] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[27][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(SyncReset_X58_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan56~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][1] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[24][1] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][1] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][1] .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|pwmList[24][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[27][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan56~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(SyncReset_X58_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan56~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][2] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[24][2] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][2] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[24][2] .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|pwmList[24][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][3] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[24][3]~q ),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan50~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X56_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y9_SIG ),
	.SyncReset(SyncReset_X56_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan50~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][3] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[24][3] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][3] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[24][3] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[24][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[24][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan50~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X56_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y9_SIG ),
	.SyncReset(SyncReset_X56_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan50~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][4] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[24][4] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][4] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[24][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[24][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X56_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[24][5]~56_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][5] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[24][5] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][5] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[24][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[24][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[24][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan50~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X56_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y9_SIG ),
	.SyncReset(SyncReset_X56_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y9_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan50~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][6] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[24][6] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][6] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[24][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[24][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][7] (
	.A(\macro_inst|controller|sm_pwm|pwmList[24][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan50~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X56_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y9_SIG ),
	.SyncReset(SyncReset_X56_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan50~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][7] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[24][7] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][7] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[24][7] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[24][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][7] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[24][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(SyncReset_X58_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan49~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][8] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[24][8] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][8] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[24][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[24][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[24][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan49~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[24][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~56_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(SyncReset_X58_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan49~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[24][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[24][9] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[24][9] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[24][9] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[24][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[24][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[24][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[24][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[25][0]~9_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][0] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][0] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[25][0] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[25][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[25][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[25][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan51~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(SyncReset_X61_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan51~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][10] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][10] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][10] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[25][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[25][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[25][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan51~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(SyncReset_X61_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan51~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][11] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][11] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][11] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[25][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[25][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[25][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan51~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(SyncReset_X61_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan51~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][12] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][12] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][12] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[25][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[25][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[25][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan51~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(SyncReset_X61_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan51~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][13] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][13] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][13] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[25][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[25][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[25][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan51~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(SyncReset_X61_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan51~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][14] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][14] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][14] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[25][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[25][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][15] (
	.A(\macro_inst|ahb_add_reg [3]),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|ahb_add_reg [2]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X60_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y3_SIG ),
	.SyncReset(SyncReset_X60_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][15] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][15] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[25][15] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[25][15] .mask = 16'h5500;
defparam \macro_inst|controller|sm_pwm|pwmList[25][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[25][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan52~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y2_SIG ),
	.SyncReset(SyncReset_X61_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan52~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][1] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][1] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[25][1] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[25][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[25][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[25][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan52~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y2_SIG ),
	.SyncReset(SyncReset_X61_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan52~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][2] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][2] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[25][2] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[25][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[25][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[25][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan52~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y2_SIG ),
	.SyncReset(SyncReset_X61_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan52~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][3] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][3] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[25][3] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[25][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[25][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[25][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan52~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y2_SIG ),
	.SyncReset(SyncReset_X61_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan52~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][4] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][4] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[25][4] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[25][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[25][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X60_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[25][5]~8_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][5] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][5] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[25][5] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[25][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[25][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[25][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan52~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y2_SIG ),
	.SyncReset(SyncReset_X61_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y2_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan52~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][6] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][6] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[25][6] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[25][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[25][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][7] (
	.A(vcc),
	.B(\macro_inst|ahb_add_reg [3]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|ahb_add_reg [2]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X60_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y3_SIG ),
	.SyncReset(SyncReset_X60_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~15_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][7] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][7] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[25][7] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[25][7] .mask = 16'h00CC;
defparam \macro_inst|controller|sm_pwm|pwmList[25][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[25][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(SyncReset_X61_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan51~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][8] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][8] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][8] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[25][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[25][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[25][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan51~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[25][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~80_combout_X61_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y3_SIG ),
	.SyncReset(SyncReset_X61_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan51~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[25][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[25][9] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[25][9] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][9] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[25][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[25][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[25][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[25][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X56_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[26][0]~59_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][0] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[26][0] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[26][0] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[26][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[26][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[26][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan53~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(SyncReset_X60_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan53~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][10] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[26][10] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[26][10] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[26][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[26][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[26][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan53~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(SyncReset_X60_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan53~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][11] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[26][11] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[26][11] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[26][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[26][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[26][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan53~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(SyncReset_X60_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan53~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][12] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[26][12] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[26][12] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[26][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[26][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[26][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan53~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(SyncReset_X60_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan53~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][13] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[26][13] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[26][13] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[26][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[26][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[26][14]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan53~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(SyncReset_X60_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y10_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan53~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][14] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[26][14] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[26][14] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[26][14] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[26][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[26][7]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X56_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ),
	.SyncReset(SyncReset_X56_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y6_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~178_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][15] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[26][15] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[26][15] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[26][15] .mask = 16'hFFD1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][1] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[26][1]~q ),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan54~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X56_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ),
	.SyncReset(SyncReset_X56_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan54~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][1] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[26][1] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[26][1] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[26][1] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[26][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][2] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.B(\macro_inst|controller|sm_pwm|pwmList[26][2]~q ),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan54~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X56_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ),
	.SyncReset(SyncReset_X56_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan54~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][2] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[26][2] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[26][2] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[26][2] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[26][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[26][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan54~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X56_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ),
	.SyncReset(SyncReset_X56_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan54~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][3] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[26][3] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[26][3] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[26][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[26][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[26][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan54~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X56_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ),
	.SyncReset(SyncReset_X56_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan54~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][4] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[26][4] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[26][4] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[26][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[26][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X56_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[26][5]~58_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][5] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[26][5] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[26][5] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[26][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[26][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[26][6]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan54~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X56_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ),
	.SyncReset(SyncReset_X56_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y6_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan54~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][6] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[26][6] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[26][6] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[26][6] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[26][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X56_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[26][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][7] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[26][7] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[26][7] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[26][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[26][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[26][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(SyncReset_X60_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan53~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][8] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[26][8] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[26][8] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[26][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[26][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[26][9] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[26][9]~q ),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan53~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[26][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~57_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(SyncReset_X60_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan53~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[26][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[26][9] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[26][9] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[26][9] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[26][9] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[26][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[26][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[26][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[27][0]~11_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][0] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[27][0] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[27][0] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[27][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][10] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[10] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[27][10]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][10] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[27][10] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[27][10] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[27][10] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[27][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][10] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][10] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][11] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[11] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[27][11]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][11] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[27][11] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[27][11] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[27][11] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[27][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][11] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][11] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][12] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[12] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[27][12]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][12] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[27][12] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[27][12] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[27][12] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[27][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][12] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][12] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][13] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[13] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[27][13]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][13] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[27][13] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[27][13] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[27][13] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[27][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][13] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][13] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][14] (
	.A(\macro_inst|controller|sm_pwm|pwmList[34][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan70~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y8_SIG ),
	.SyncReset(SyncReset_X58_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan70~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][14] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[27][14] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[27][14] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[27][14] .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|pwmList[27][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][14] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][15] (
	.A(\macro_inst|controller|sm_pwm|LessThan56~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[27][7]~q ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X57_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y8_SIG ),
	.SyncReset(SyncReset_X57_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y8_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~82_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][15] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[27][15] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[27][15] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[27][15] .mask = 16'h77F0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[27][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan56~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(SyncReset_X58_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan56~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][1] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[27][1] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[27][1] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[27][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[27][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[27][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan56~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(SyncReset_X58_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan56~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][2] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[27][2] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[27][2] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[27][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[27][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[27][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan56~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(SyncReset_X58_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan56~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][3] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[27][3] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[27][3] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[27][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[27][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[27][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan56~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(SyncReset_X58_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan56~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][4] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[27][4] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[27][4] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[27][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[27][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[27][5]~10_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][5] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[27][5] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[27][5] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[27][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[27][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[27][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan56~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y9_SIG ),
	.SyncReset(SyncReset_X58_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y9_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan56~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][6] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[27][6] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[27][6] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[27][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[27][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][7] (
	.A(\macro_inst|ahb_add_reg [1]),
	.B(\macro_inst|ahb_add_reg [4]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|ahb_add_reg [5]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X58_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y8_SIG ),
	.SyncReset(SyncReset_X58_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y8_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~22_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][7] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[27][7] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[27][7] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[27][7] .mask = 16'h8800;
defparam \macro_inst|controller|sm_pwm|pwmList[27][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[27][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X57_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y8_SIG ),
	.SyncReset(SyncReset_X57_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan55~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][8] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[27][8] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[27][8] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[27][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[27][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[27][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan55~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[27][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~23_combout_X57_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y8_SIG ),
	.SyncReset(SyncReset_X57_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan55~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[27][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[27][9] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[27][9] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[27][9] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[27][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[27][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[27][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[28][0]~61_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][0] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[28][0] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[28][0] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[28][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[28][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][10] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.B(\macro_inst|controller|sm_pwm|pwmList[28][10]~q ),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan57~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ),
	.SyncReset(SyncReset_X56_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan57~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][10] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[28][10] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][10] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[28][10] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[28][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[28][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan57~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ),
	.SyncReset(SyncReset_X56_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan57~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][11] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[28][11] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][11] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[28][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[28][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[28][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan57~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ),
	.SyncReset(SyncReset_X56_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan57~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][12] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[28][12] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][12] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[28][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[28][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[28][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan57~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ),
	.SyncReset(SyncReset_X56_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan57~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][13] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[28][13] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][13] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[28][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[28][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[28][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan57~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ),
	.SyncReset(SyncReset_X56_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y8_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan57~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][14] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[28][14] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][14] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[28][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[28][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[28][7]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|LessThan58~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ),
	.SyncReset(SyncReset_X56_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~228_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][15] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[28][15] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[28][15] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[28][15] .mask = 16'h74FC;
defparam \macro_inst|controller|sm_pwm|pwmList[28][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[28][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan58~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ),
	.SyncReset(SyncReset_X56_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan58~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][1] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[28][1] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[28][1] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[28][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[28][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][2] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.B(\macro_inst|controller|sm_pwm|pwmList[28][2]~q ),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan58~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ),
	.SyncReset(SyncReset_X56_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan58~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][2] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[28][2] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[28][2] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[28][2] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[28][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[28][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan58~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ),
	.SyncReset(SyncReset_X56_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan58~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][3] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[28][3] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[28][3] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[28][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[28][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[28][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan58~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ),
	.SyncReset(SyncReset_X56_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan58~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][4] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[28][4] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[28][4] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[28][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[28][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[28][5]~60_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][5] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[28][5] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[28][5] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[28][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[28][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[28][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan58~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ),
	.SyncReset(SyncReset_X56_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan58~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][6] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[28][6] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[28][6] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[28][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[28][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][7] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[28][15]~q ),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|LessThan57~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y7_SIG ),
	.SyncReset(SyncReset_X56_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~180_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][7] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[28][7] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[28][7] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[28][7] .mask = 16'h8DAF;
defparam \macro_inst|controller|sm_pwm|pwmList[28][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[28][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ),
	.SyncReset(SyncReset_X56_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan57~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][8] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[28][8] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][8] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[28][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[28][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[28][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[28][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan57~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[28][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~58_combout_X56_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ),
	.SyncReset(SyncReset_X56_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan57~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[28][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[28][9] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[28][9] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][9] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[28][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[28][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[28][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[28][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][0] (
	.A(\rv32.mem_ahb_hwdata[0] ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X58_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[29][0]~13_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][0] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[29][0] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[29][0] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[29][0] .mask = 16'h5555;
defparam \macro_inst|controller|sm_pwm|pwmList[29][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[29][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan59~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X60_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ),
	.SyncReset(SyncReset_X60_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan59~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][10] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[29][10] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[29][10] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[29][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[29][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[29][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan59~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X60_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ),
	.SyncReset(SyncReset_X60_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan59~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][11] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[29][11] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[29][11] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[29][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[29][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][12] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[29][12]~q ),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan59~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X60_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ),
	.SyncReset(SyncReset_X60_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan59~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][12] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[29][12] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[29][12] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[29][12] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[29][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[29][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan59~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X60_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ),
	.SyncReset(SyncReset_X60_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan59~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][13] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[29][13] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[29][13] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[29][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[29][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[29][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan59~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X60_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ),
	.SyncReset(SyncReset_X60_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y5_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan59~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][14] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[29][14] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[29][14] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[29][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[29][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][15] (
	.A(\macro_inst|controller|sm_pwm|LessThan60~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[29][7]~q ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X58_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y5_SIG ),
	.SyncReset(SyncReset_X58_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y5_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~84_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][15] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[29][15] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[29][15] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[29][15] .mask = 16'h77F0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][1] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[29][1]~q ),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan60~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X58_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y5_SIG ),
	.SyncReset(SyncReset_X58_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan60~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][1] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[29][1] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[29][1] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][1] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[29][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[29][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan60~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X58_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y5_SIG ),
	.SyncReset(SyncReset_X58_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan60~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][2] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[29][2] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[29][2] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[29][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[29][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][3] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[29][3]~q ),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan60~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X58_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y5_SIG ),
	.SyncReset(SyncReset_X58_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan60~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][3] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[29][3] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[29][3] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[29][3] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[29][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][4] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X58_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y5_SIG ),
	.SyncReset(SyncReset_X58_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y5_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[4]~4_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][4] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[29][4] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[29][4] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[29][4] .mask = 16'hCC00;
defparam \macro_inst|controller|sm_pwm|pwmList[29][4] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][4] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][5] (
	.A(vcc),
	.B(\rv32.mem_ahb_hwdata[5] ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X58_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[29][5]~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][5] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[29][5] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[29][5] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[29][5] .mask = 16'h3333;
defparam \macro_inst|controller|sm_pwm|pwmList[29][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][6] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [6]),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X58_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y5_SIG ),
	.SyncReset(SyncReset_X58_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y5_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[6]~6_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][6] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[29][6] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[29][6] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[29][6] .mask = 16'hCC00;
defparam \macro_inst|controller|sm_pwm|pwmList[29][6] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][7] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [7]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X58_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y5_SIG ),
	.SyncReset(SyncReset_X58_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y5_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[7]~7_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][7] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[29][7] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[29][7] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[29][7] .mask = 16'hCC00;
defparam \macro_inst|controller|sm_pwm|pwmList[29][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[29][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X60_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ),
	.SyncReset(SyncReset_X60_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan59~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][8] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[29][8] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[29][8] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[29][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[29][9] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[29][9]~q ),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan59~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[29][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~24_combout_X60_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ),
	.SyncReset(SyncReset_X60_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan59~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[29][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[29][9] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[29][9] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[29][9] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][9] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[29][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[29][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[29][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X56_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[2][0]~51_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][0] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[2][0] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][0] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[2][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][10] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.B(\macro_inst|controller|sm_pwm|pwmList[2][2]~q ),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan6~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X56_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ),
	.SyncReset(SyncReset_X56_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan6~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][10] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[2][10] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][10] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[2][10] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[2][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[2][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan5~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(SyncReset_X57_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan5~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][11] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[2][11] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][11] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[2][11] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[2][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][12] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[12] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X56_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[2][12]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][12] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[2][12] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][12] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[2][12] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[2][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][12] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][12] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][13] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[2][11]~q ),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan5~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(SyncReset_X57_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan5~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][13] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[2][13] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][13] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[2][13] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[2][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][14] (
	.A(\macro_inst|controller|sm_pwm|pwmList[2][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan6~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X56_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ),
	.SyncReset(SyncReset_X56_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan6~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][14] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[2][14] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][14] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[2][14] .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|pwmList[2][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][14] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[2][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan5~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(SyncReset_X57_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan5~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][15] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[2][15] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][15] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[2][15] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[2][15] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][15] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][1] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[2][9]~q ),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan5~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(SyncReset_X57_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan5~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][1] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[2][1] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][1] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[2][1] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[2][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][2] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[2][14]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan5~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(SyncReset_X57_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y10_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan5~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][2] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[2][2] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][2] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[2][2] .mask = 16'h5F05;
defparam \macro_inst|controller|sm_pwm|pwmList[2][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][2] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[2][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan6~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X56_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ),
	.SyncReset(SyncReset_X56_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan6~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][3] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[2][3] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][3] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[2][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[2][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[2][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan6~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X56_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ),
	.SyncReset(SyncReset_X56_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan6~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][4] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[2][4] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][4] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[2][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[2][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X56_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[2][5]~50_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][5] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[2][5] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][5] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[2][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[2][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[2][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan6~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X56_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ),
	.SyncReset(SyncReset_X56_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y10_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan6~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][6] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[2][6] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][6] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[2][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[2][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][7] (
	.A(\macro_inst|controller|sm_pwm|pwmList[2][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan6~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X56_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y10_SIG ),
	.SyncReset(SyncReset_X56_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan6~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][7] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[2][7] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][7] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[2][7] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[2][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][7] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[2][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(SyncReset_X57_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan5~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][8] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[2][8] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][8] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[2][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[2][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[2][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[2][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan5~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[2][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~50_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(SyncReset_X57_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan5~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[2][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[2][9] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[2][9] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[2][9] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[2][9] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[2][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[2][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[2][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X57_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[30][0]~63_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][0] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[30][0] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[30][0] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[30][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[30][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[30][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan61~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X60_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ),
	.SyncReset(SyncReset_X60_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan61~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][10] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[30][10] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[30][10] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[30][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[30][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[30][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan61~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X60_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ),
	.SyncReset(SyncReset_X60_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan61~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][11] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[30][11] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[30][11] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[30][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[30][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][12] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[30][12]~q ),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan61~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X60_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ),
	.SyncReset(SyncReset_X60_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan61~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][12] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[30][12] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[30][12] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[30][12] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[30][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[30][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan61~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X60_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ),
	.SyncReset(SyncReset_X60_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan61~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][13] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[30][13] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[30][13] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[30][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[30][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[30][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan61~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X60_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ),
	.SyncReset(SyncReset_X60_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y5_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan61~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][14] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[30][14] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[30][14] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[30][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[30][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[30][7]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan62~12_combout ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X57_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ),
	.SyncReset(SyncReset_X57_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y9_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~230_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][15] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[30][15] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[30][15] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[30][15] .mask = 16'h77F0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[30][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan62~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X57_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ),
	.SyncReset(SyncReset_X57_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan62~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][1] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[30][1] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[30][1] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[30][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[30][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan62~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X57_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ),
	.SyncReset(SyncReset_X57_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan62~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][2] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[30][2] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[30][2] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[30][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[30][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[30][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan62~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X57_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ),
	.SyncReset(SyncReset_X57_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan62~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][3] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[30][3] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[30][3] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[30][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[30][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[30][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan62~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X57_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ),
	.SyncReset(SyncReset_X57_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan62~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][4] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[30][4] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[30][4] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[30][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[30][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][5] (
	.A(\rv32.mem_ahb_hwdata[5] ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X57_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[30][5]~62_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][5] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[30][5] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[30][5] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[30][5] .mask = 16'h5555;
defparam \macro_inst|controller|sm_pwm|pwmList[30][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[30][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan62~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X57_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ),
	.SyncReset(SyncReset_X57_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y9_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan62~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][6] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[30][6] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[30][6] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[30][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[30][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X57_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[30][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][7] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[30][7] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[30][7] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[30][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[30][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[30][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X60_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ),
	.SyncReset(SyncReset_X60_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan61~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][8] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[30][8] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[30][8] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[30][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[30][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[30][9] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[30][9]~q ),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan61~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[30][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~59_combout_X60_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y5_SIG ),
	.SyncReset(SyncReset_X60_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan61~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[30][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[30][9] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[30][9] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[30][9] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[30][9] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[30][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[30][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[30][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[31][0]~15_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][0] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[31][0] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][0] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[31][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[31][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan63~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X57_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ),
	.SyncReset(SyncReset_X57_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan63~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][10] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[31][10] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][10] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[31][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[31][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[31][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan63~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X57_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ),
	.SyncReset(SyncReset_X57_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan63~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][11] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[31][11] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][11] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[31][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[31][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][12] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[31][12]~q ),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan63~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X57_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ),
	.SyncReset(SyncReset_X57_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan63~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][12] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[31][12] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][12] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[31][12] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[31][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[31][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan63~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X57_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ),
	.SyncReset(SyncReset_X57_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan63~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][13] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[31][13] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][13] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[31][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[31][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[31][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan63~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X57_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ),
	.SyncReset(SyncReset_X57_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y11_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan63~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][14] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[31][14] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][14] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[31][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[31][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[31][7]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan64~12_combout ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X57_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ),
	.SyncReset(SyncReset_X57_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y11_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~86_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][15] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[31][15] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][15] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[31][15] .mask = 16'h77F0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[31][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan64~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(SyncReset_X59_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan64~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][1] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[31][1] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][1] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[31][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[31][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan64~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(SyncReset_X59_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan64~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][2] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[31][2] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][2] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[31][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[31][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[31][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan64~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(SyncReset_X59_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan64~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][3] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[31][3] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][3] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[31][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[31][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[31][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan64~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(SyncReset_X59_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan64~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][4] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[31][4] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][4] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[31][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[31][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[31][5]~14_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][5] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[31][5] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][5] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[31][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[31][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan64~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X59_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y9_SIG ),
	.SyncReset(SyncReset_X59_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y9_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan64~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][6] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[31][6] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][6] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[31][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[31][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][7] (
	.A(\macro_inst|controller|sm_pwm|pwmList[31][15]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan63~12_combout ),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X57_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ),
	.SyncReset(SyncReset_X57_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y11_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~38_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][7] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[31][7] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][7] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][7] .mask = 16'hBB0F;
defparam \macro_inst|controller|sm_pwm|pwmList[31][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[31][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X57_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ),
	.SyncReset(SyncReset_X57_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan63~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][8] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[31][8] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][8] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[31][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[31][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[31][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[31][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan63~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[31][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~25_combout_X57_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y11_SIG ),
	.SyncReset(SyncReset_X57_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan63~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[31][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[31][9] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[31][9] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][9] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[31][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[31][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[31][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[31][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[32][0]~65_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][0] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[32][0] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[32][0] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[32][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[32][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[32][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan65~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(SyncReset_X60_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan65~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][10] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[32][10] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[32][10] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[32][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[32][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[32][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan65~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(SyncReset_X60_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan65~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][11] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[32][11] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[32][11] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[32][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[32][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[32][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan65~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(SyncReset_X60_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan65~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][12] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[32][12] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[32][12] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[32][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[32][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[32][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan65~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(SyncReset_X60_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan65~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][13] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[32][13] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[32][13] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[32][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[32][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[32][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan65~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(SyncReset_X60_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y9_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan65~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][14] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[32][14] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[32][14] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[32][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[32][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][15] (
	.A(\macro_inst|controller|sm_pwm|LessThan66~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[32][7]~q ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X61_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ),
	.SyncReset(SyncReset_X61_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y9_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~232_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][15] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[32][15] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[32][15] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[32][15] .mask = 16'h77F0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[32][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan66~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X61_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ),
	.SyncReset(SyncReset_X61_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan66~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][1] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[32][1] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[32][1] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[32][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[32][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[32][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan66~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X61_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ),
	.SyncReset(SyncReset_X61_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan66~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][2] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[32][2] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[32][2] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[32][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[32][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[32][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan66~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X61_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ),
	.SyncReset(SyncReset_X61_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan66~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][3] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[32][3] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[32][3] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[32][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[32][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[32][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan66~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X61_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ),
	.SyncReset(SyncReset_X61_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan66~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][4] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[32][4] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[32][4] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[32][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[32][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X61_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[32][5]~64_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][5] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[32][5] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[32][5] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[32][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[32][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[32][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan66~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X61_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ),
	.SyncReset(SyncReset_X61_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y9_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan66~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][6] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[32][6] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[32][6] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[32][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[32][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][7] (
	.A(\macro_inst|controller|sm_pwm|LessThan65~12_combout ),
	.B(\macro_inst|controller|sm_pwm|pwmList[32][15]~q ),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X61_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y9_SIG ),
	.SyncReset(SyncReset_X61_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y9_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~184_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][7] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[32][7] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[32][7] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[32][7] .mask = 16'hDD0F;
defparam \macro_inst|controller|sm_pwm|pwmList[32][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[32][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(SyncReset_X60_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan65~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][8] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[32][8] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[32][8] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[32][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[32][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[32][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[32][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan65~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[32][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~60_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(SyncReset_X60_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan65~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[32][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[32][9] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[32][9] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[32][9] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[32][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[32][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[32][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[32][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X59_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[33][0]~17_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][0] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][0] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[33][0] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[33][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[33][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[33][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan67~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X60_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ),
	.SyncReset(SyncReset_X60_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan67~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][10] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][10] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[33][10] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[33][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[33][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[33][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan67~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X60_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ),
	.SyncReset(SyncReset_X60_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan67~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][11] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][11] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[33][11] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[33][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[33][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][12] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[33][5]~q ),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan68~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X59_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ),
	.SyncReset(SyncReset_X59_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan68~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][12] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][12] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[33][12] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[33][12] .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|pwmList[33][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[33][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan67~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X60_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ),
	.SyncReset(SyncReset_X60_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan67~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][13] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][13] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[33][13] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[33][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[33][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[33][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan67~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X60_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ),
	.SyncReset(SyncReset_X60_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y12_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan67~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][14] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][14] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[33][14] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[33][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[33][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[33][7]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|LessThan68~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X59_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ),
	.SyncReset(SyncReset_X59_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y12_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~88_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][15] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][15] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[33][15] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[33][15] .mask = 16'h74FC;
defparam \macro_inst|controller|sm_pwm|pwmList[33][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[33][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan68~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X59_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ),
	.SyncReset(SyncReset_X59_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan68~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][1] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][1] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[33][1] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[33][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[33][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan68~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X59_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ),
	.SyncReset(SyncReset_X59_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan68~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][2] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][2] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[33][2] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[33][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[33][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][3] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[33][3]~q ),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan68~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X59_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ),
	.SyncReset(SyncReset_X59_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan68~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][3] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][3] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[33][3] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[33][3] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[33][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[33][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan68~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X59_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ),
	.SyncReset(SyncReset_X59_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan68~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][4] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][4] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[33][4] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[33][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[33][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X59_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[33][5]~16_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][5] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][5] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[33][5] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[33][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[33][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[33][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan68~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X59_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ),
	.SyncReset(SyncReset_X59_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y12_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan68~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][6] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][6] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[33][6] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[33][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[33][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][7] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[33][15]~q ),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|LessThan67~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X59_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y12_SIG ),
	.SyncReset(SyncReset_X59_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y12_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~40_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][7] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][7] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[33][7] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[33][7] .mask = 16'h8DAF;
defparam \macro_inst|controller|sm_pwm|pwmList[33][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][8] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[8] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X60_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[33][8]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][8] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][8] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[33][8] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[33][8] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[33][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][8] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][8] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[33][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[33][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan67~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[33][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~28_combout_X60_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ),
	.SyncReset(SyncReset_X60_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan67~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[33][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[33][9] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[33][9] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[33][9] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[33][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[33][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[33][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][0] (
	.A(\rv32.mem_ahb_hwdata[0] ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X56_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[34][0]~67_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][0] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[34][0] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[34][0] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[34][0] .mask = 16'h5555;
defparam \macro_inst|controller|sm_pwm|pwmList[34][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[34][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan69~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X56_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ),
	.SyncReset(SyncReset_X56_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan69~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][10] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[34][10] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[34][10] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[34][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[34][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[34][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan69~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X56_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ),
	.SyncReset(SyncReset_X56_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan69~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][11] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[34][11] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[34][11] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[34][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[34][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][12] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[12] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X56_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[34][12]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][12] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[34][12] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[34][12] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[34][12] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[34][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][12] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][12] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[34][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan69~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X56_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ),
	.SyncReset(SyncReset_X56_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan69~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][13] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[34][13] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[34][13] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[34][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[34][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[34][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan69~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X56_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ),
	.SyncReset(SyncReset_X56_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan69~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][14] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[34][14] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[34][14] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[34][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[34][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[1][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan4~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X59_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ),
	.SyncReset(SyncReset_X59_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan4~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][15] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[34][15] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[34][15] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[34][15] .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|pwmList[34][15] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][15] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][1] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[1] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X59_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[34][1]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][1] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[34][1] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[34][1] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][1] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[34][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][1] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][1] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][2] (
	.A(\macro_inst|ahb_add_reg [5]),
	.B(\macro_inst|ahb_add_reg [6]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(\macro_inst|ahb_add_reg [4]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X59_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ),
	.SyncReset(SyncReset_X59_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~32_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][2] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[34][2] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[34][2] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][2] .mask = 16'h0044;
defparam \macro_inst|controller|sm_pwm|pwmList[34][2] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][2] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][3] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[3] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X59_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[34][3]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][3] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[34][3] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[34][3] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[34][3] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[34][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][3] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][3] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][4] (
	.A(\macro_inst|ahb_add_reg [5]),
	.B(\macro_inst|ahb_add_reg [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(\macro_inst|ahb_add_reg [6]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X59_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ),
	.SyncReset(SyncReset_X59_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~41_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][4] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[34][4] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[34][4] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[34][4] .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|pwmList[34][4] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][4] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X56_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[34][5]~66_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][5] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[34][5] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[34][5] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[34][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[34][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][6] (
	.A(\macro_inst|ahb_add_reg [5]),
	.B(\macro_inst|ahb_add_reg [4]),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|ahb_add_reg [1]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X59_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ),
	.SyncReset(SyncReset_X59_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~19_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][6] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[34][6] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[34][6] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[34][6] .mask = 16'h2200;
defparam \macro_inst|controller|sm_pwm|pwmList[34][6] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][7] (
	.A(\macro_inst|controller|sm_pwm|pwmList[1][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X59_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y7_SIG ),
	.SyncReset(SyncReset_X59_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan4~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][7] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[34][7] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[34][7] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[34][7] .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|pwmList[34][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][7] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[34][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X56_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ),
	.SyncReset(SyncReset_X56_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan69~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][8] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[34][8] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[34][8] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[34][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[34][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[34][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[34][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan69~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[34][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~61_combout_X56_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y4_SIG ),
	.SyncReset(SyncReset_X56_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan69~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[34][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[34][9] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[34][9] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[34][9] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[34][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[34][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[34][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[34][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X58_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[35][0]~19_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][0] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][0] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[35][0] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[35][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[35][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[35][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan71~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X57_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(SyncReset_X57_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan71~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][10] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][10] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[35][10] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[35][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[35][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[35][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan71~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X57_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(SyncReset_X57_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan71~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][11] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][11] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[35][11] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[35][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[35][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][12] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[35][12]~q ),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan71~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X57_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(SyncReset_X57_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan71~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][12] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][12] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[35][12] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[35][12] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[35][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][13] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[35][13]~q ),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan71~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X57_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(SyncReset_X57_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan71~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][13] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][13] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[35][13] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[35][13] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[35][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[35][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan71~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X57_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(SyncReset_X57_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan71~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][14] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][14] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[35][14] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[35][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[35][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][15] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[15] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X57_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[35][15]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][15] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][15] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[35][15] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[35][15] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[35][15] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][15] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[35][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan72~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X58_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ),
	.SyncReset(SyncReset_X58_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan72~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][1] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][1] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[35][1] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[35][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[35][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[35][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan72~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X58_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ),
	.SyncReset(SyncReset_X58_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan72~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][2] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][2] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[35][2] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[35][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[35][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[35][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan72~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X58_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ),
	.SyncReset(SyncReset_X58_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan72~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][3] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][3] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[35][3] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[35][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[35][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[35][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan72~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X58_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ),
	.SyncReset(SyncReset_X58_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan72~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][4] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][4] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[35][4] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[35][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[35][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X58_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[35][5]~18_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][5] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][5] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[35][5] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[35][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[35][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[35][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan72~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X58_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ),
	.SyncReset(SyncReset_X58_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y2_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan72~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][6] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][6] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[35][6] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[35][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[35][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][7] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[35][15]~q ),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|LessThan71~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X57_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(SyncReset_X57_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~42_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][7] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][7] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[35][7] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[35][7] .mask = 16'h8DAF;
defparam \macro_inst|controller|sm_pwm|pwmList[35][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][8] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[35][8]~q ),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X57_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(SyncReset_X57_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan71~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][8] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][8] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[35][8] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][8] .mask = 16'h0044;
defparam \macro_inst|controller|sm_pwm|pwmList[35][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[35][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[35][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan71~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[35][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~30_combout_X57_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y4_SIG ),
	.SyncReset(SyncReset_X57_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan71~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[35][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[35][9] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[35][9] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[35][9] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[35][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[35][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[35][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[35][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X58_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[36][0]~69_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][0] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[36][0] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[36][0] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[36][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[36][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[36][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan73~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X57_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y8_SIG ),
	.SyncReset(SyncReset_X57_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan73~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][10] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[36][10] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[36][10] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[36][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[36][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[36][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan73~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X57_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y8_SIG ),
	.SyncReset(SyncReset_X57_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan73~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][11] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[36][11] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[36][11] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[36][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[36][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][12] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[36][12]~q ),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan73~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X57_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y8_SIG ),
	.SyncReset(SyncReset_X57_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan73~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][12] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[36][12] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[36][12] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[36][12] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[36][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[36][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan73~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X57_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y8_SIG ),
	.SyncReset(SyncReset_X57_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan73~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][13] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[36][13] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[36][13] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[36][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[36][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[36][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan73~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X57_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y8_SIG ),
	.SyncReset(SyncReset_X57_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y8_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan73~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][14] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[36][14] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[36][14] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[36][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[36][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][15] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[36][7]~q ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|LessThan74~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X58_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y7_SIG ),
	.SyncReset(SyncReset_X58_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~236_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][15] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[36][15] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[36][15] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[36][15] .mask = 16'h72FA;
defparam \macro_inst|controller|sm_pwm|pwmList[36][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][1] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[36][1]~q ),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan74~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X58_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y7_SIG ),
	.SyncReset(SyncReset_X58_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan74~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][1] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[36][1] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[36][1] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][1] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[36][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[36][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan74~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X58_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y7_SIG ),
	.SyncReset(SyncReset_X58_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan74~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][2] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[36][2] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[36][2] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[36][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[36][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[36][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan74~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X58_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y7_SIG ),
	.SyncReset(SyncReset_X58_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan74~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][3] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[36][3] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[36][3] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[36][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[36][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[36][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan74~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X58_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y7_SIG ),
	.SyncReset(SyncReset_X58_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan74~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][4] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[36][4] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[36][4] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[36][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[36][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X58_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[36][5]~68_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][5] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[36][5] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[36][5] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[36][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[36][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[36][6]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan74~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X58_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y7_SIG ),
	.SyncReset(SyncReset_X58_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan74~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][6] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[36][6] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[36][6] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[36][6] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[36][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][7] (
	.A(\macro_inst|controller|sm_pwm|pwmList[36][15]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|LessThan73~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X58_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y7_SIG ),
	.SyncReset(SyncReset_X58_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~188_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][7] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[36][7] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[36][7] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[36][7] .mask = 16'h8BCF;
defparam \macro_inst|controller|sm_pwm|pwmList[36][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[36][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X57_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y8_SIG ),
	.SyncReset(SyncReset_X57_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan73~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][8] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[36][8] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[36][8] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[36][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[36][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[36][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[36][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan73~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[36][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~62_combout_X57_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y8_SIG ),
	.SyncReset(SyncReset_X57_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan73~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[36][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[36][9] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[36][9] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[36][9] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[36][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[36][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[36][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[36][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][0] (
	.A(vcc),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[0] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X61_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[37][0]~21_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][0] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[37][0] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][0] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[37][0] .mask = 16'h0F0F;
defparam \macro_inst|controller|sm_pwm|pwmList[37][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[37][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan75~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(SyncReset_X60_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan75~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][10] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[37][10] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[37][10] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[37][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[37][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[37][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan75~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(SyncReset_X60_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan75~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][11] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[37][11] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[37][11] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[37][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[37][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[37][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan75~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(SyncReset_X60_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan75~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][12] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[37][12] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[37][12] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[37][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[37][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[37][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan75~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(SyncReset_X60_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan75~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][13] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[37][13] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[37][13] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[37][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[37][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[37][14]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan75~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(SyncReset_X60_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y2_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan75~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][14] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[37][14] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[37][14] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[37][14] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[37][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][15] (
	.A(\macro_inst|controller|sm_pwm|LessThan76~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[37][7]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X61_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ),
	.SyncReset(SyncReset_X61_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y5_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~92_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][15] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[37][15] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][15] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[37][15] .mask = 16'h74FC;
defparam \macro_inst|controller|sm_pwm|pwmList[37][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[37][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan76~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X61_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ),
	.SyncReset(SyncReset_X61_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan76~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][1] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[37][1] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][1] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[37][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[37][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan76~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X61_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ),
	.SyncReset(SyncReset_X61_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan76~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][2] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[37][2] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][2] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[37][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[37][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[37][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan76~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X61_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ),
	.SyncReset(SyncReset_X61_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan76~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][3] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[37][3] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][3] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[37][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[37][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[37][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan76~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X61_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ),
	.SyncReset(SyncReset_X61_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan76~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][4] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[37][4] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][4] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[37][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[37][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X61_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[37][5]~20_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][5] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[37][5] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][5] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[37][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[37][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[37][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan76~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X61_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ),
	.SyncReset(SyncReset_X61_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y5_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan76~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][6] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[37][6] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][6] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[37][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[37][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X61_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[37][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][7] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[37][7] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][7] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[37][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[37][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[37][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(SyncReset_X60_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan75~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][8] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[37][8] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[37][8] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[37][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[37][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[37][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[37][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan75~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[37][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~31_combout_X60_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y2_SIG ),
	.SyncReset(SyncReset_X60_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan75~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[37][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[37][9] .coord_x = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[37][9] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[37][9] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[37][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[37][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[37][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[37][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][0] (
	.A(vcc),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[0] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[38][0]~71_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][0] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[38][0] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[38][0] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[38][0] .mask = 16'h0F0F;
defparam \macro_inst|controller|sm_pwm|pwmList[38][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[38][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan77~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan77~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][10] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[38][10] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[38][10] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[38][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[38][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][11] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[38][11]~q ),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan77~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan77~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][11] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[38][11] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[38][11] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[38][11] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[38][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[38][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan77~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan77~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][12] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[38][12] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[38][12] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[38][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[38][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[38][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan77~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan77~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][13] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[38][13] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[38][13] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[38][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[38][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[38][14]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan77~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan77~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][14] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[38][14] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[38][14] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[38][14] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[38][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[38][7]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|LessThan78~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X62_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ),
	.SyncReset(SyncReset_X62_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y5_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~238_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][15] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[38][15] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[38][15] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[38][15] .mask = 16'h74FC;
defparam \macro_inst|controller|sm_pwm|pwmList[38][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[38][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan78~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X62_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ),
	.SyncReset(SyncReset_X62_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan78~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][1] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[38][1] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[38][1] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[38][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[38][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[38][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan78~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X62_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ),
	.SyncReset(SyncReset_X62_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan78~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][2] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[38][2] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[38][2] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[38][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[38][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[38][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan78~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X62_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ),
	.SyncReset(SyncReset_X62_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan78~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][3] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[38][3] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[38][3] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[38][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[38][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[38][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan78~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X62_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ),
	.SyncReset(SyncReset_X62_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan78~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][4] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[38][4] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[38][4] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[38][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[38][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X62_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[38][5]~70_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][5] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[38][5] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[38][5] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[38][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[38][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][6] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.B(\macro_inst|controller|sm_pwm|pwmList[38][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan78~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X62_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ),
	.SyncReset(SyncReset_X62_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y5_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan78~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][6] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[38][6] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[38][6] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[38][6] .mask = 16'h4D4D;
defparam \macro_inst|controller|sm_pwm|pwmList[38][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X62_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[38][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][7] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[38][7] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[38][7] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[38][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[38][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[38][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan77~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][8] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[38][8] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[38][8] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[38][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[38][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[38][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan77~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[38][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~64_combout_X61_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y6_SIG ),
	.SyncReset(SyncReset_X61_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan77~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[38][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[38][9] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[38][9] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[38][9] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[38][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[38][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[38][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X62_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[39][0]~23_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][0] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[39][0] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[39][0] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[39][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[39][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][10] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.B(\macro_inst|controller|sm_pwm|pwmList[39][10]~q ),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan79~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X56_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ),
	.SyncReset(SyncReset_X56_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan79~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][10] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[39][10] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][10] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[39][10] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[39][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[39][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan79~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X56_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ),
	.SyncReset(SyncReset_X56_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan79~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][11] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[39][11] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][11] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[39][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[39][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[39][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan79~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X56_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ),
	.SyncReset(SyncReset_X56_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan79~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][12] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[39][12] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][12] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[39][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[39][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[39][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan79~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X56_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ),
	.SyncReset(SyncReset_X56_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan79~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][13] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[39][13] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][13] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[39][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[39][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[39][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan79~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X56_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ),
	.SyncReset(SyncReset_X56_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y8_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan79~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][14] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[39][14] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][14] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[39][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[39][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][15] (
	.A(\macro_inst|controller|sm_pwm|LessThan80~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[39][7]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X62_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ),
	.SyncReset(SyncReset_X62_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y8_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~94_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][15] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[39][15] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[39][15] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[39][15] .mask = 16'h74FC;
defparam \macro_inst|controller|sm_pwm|pwmList[39][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[39][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan80~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X62_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ),
	.SyncReset(SyncReset_X62_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan80~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][1] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[39][1] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[39][1] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[39][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[39][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[39][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan80~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X62_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ),
	.SyncReset(SyncReset_X62_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan80~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][2] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[39][2] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[39][2] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[39][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[39][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[39][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan80~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X62_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ),
	.SyncReset(SyncReset_X62_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan80~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][3] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[39][3] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[39][3] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[39][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[39][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[39][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan80~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X62_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ),
	.SyncReset(SyncReset_X62_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan80~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][4] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[39][4] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[39][4] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[39][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[39][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X62_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[39][5]~22_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][5] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[39][5] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[39][5] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[39][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][6] (
	.A(\macro_inst|controller|sm_pwm|pwmList[39][6]~q ),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan80~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X62_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ),
	.SyncReset(SyncReset_X62_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y8_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan80~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][6] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[39][6] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[39][6] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[39][6] .mask = 16'h0AAF;
defparam \macro_inst|controller|sm_pwm|pwmList[39][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X62_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[39][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][7] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[39][7] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[39][7] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[39][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[39][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X56_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ),
	.SyncReset(SyncReset_X56_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan79~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][8] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[39][8] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][8] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[39][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[39][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[39][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[39][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan79~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[39][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~33_combout_X56_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y8_SIG ),
	.SyncReset(SyncReset_X56_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan79~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[39][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[39][9] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[39][9] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][9] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[39][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[39][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[39][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[39][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X58_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[3][0]~3_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][0] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[3][0] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[3][0] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[3][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[3][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][10] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[10] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X59_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[3][10]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][10] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[3][10] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[3][10] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[3][10] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[3][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][10] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][10] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][11] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [11]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X57_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y6_SIG ),
	.SyncReset(SyncReset_X57_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y6_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[11]~11_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][11] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[3][11] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[3][11] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[3][11] .mask = 16'hCC00;
defparam \macro_inst|controller|sm_pwm|pwmList[3][11] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][11] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[3][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan7~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X57_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y6_SIG ),
	.SyncReset(SyncReset_X57_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan7~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][12] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[3][12] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[3][12] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[3][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[3][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][13] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[13] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X59_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[3][13]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][13] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[3][13] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[3][13] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[3][13] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[3][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][13] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][13] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][14] (
	.A(\macro_inst|ahb_add_reg [6]),
	.B(\macro_inst|ahb_add_reg [5]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|ahb_add_reg [1]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X59_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y4_SIG ),
	.SyncReset(SyncReset_X59_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|Decoder0~63_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][14] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[3][14] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[3][14] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[3][14] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[3][14] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][15] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [15]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X58_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y5_SIG ),
	.SyncReset(SyncReset_X58_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y5_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[15]~15_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][15] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[3][15] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[3][15] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[3][15] .mask = 16'hCC00;
defparam \macro_inst|controller|sm_pwm|pwmList[3][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][1] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[3][1]~q ),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan8~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X58_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y3_SIG ),
	.SyncReset(SyncReset_X58_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan8~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][1] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[3][1] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[3][1] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[3][1] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[3][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[3][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan8~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X58_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y3_SIG ),
	.SyncReset(SyncReset_X58_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan8~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][2] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[3][2] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[3][2] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[3][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[3][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][3] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[3][3]~q ),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan8~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X58_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y3_SIG ),
	.SyncReset(SyncReset_X58_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan8~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][3] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[3][3] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[3][3] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[3][3] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[3][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[3][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan8~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X58_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y3_SIG ),
	.SyncReset(SyncReset_X58_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y3_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan8~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][4] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[3][4] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[3][4] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[3][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[3][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X58_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[3][5]~2_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][5] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[3][5] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[3][5] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[3][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[3][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[3][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan8~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X58_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y3_SIG ),
	.SyncReset(SyncReset_X58_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y3_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan8~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][6] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[3][6] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[3][6] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[3][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[3][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][7] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [2]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X58_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y5_SIG ),
	.SyncReset(SyncReset_X58_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y5_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[2]~2_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][7] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[3][7] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[3][7] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[3][7] .mask = 16'hCC00;
defparam \macro_inst|controller|sm_pwm|pwmList[3][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[3][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X57_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y6_SIG ),
	.SyncReset(SyncReset_X57_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan7~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][8] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[3][8] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[3][8] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[3][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[3][9] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [9]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[3][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~14_combout_X57_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y6_SIG ),
	.SyncReset(SyncReset_X57_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y6_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[9]~9_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[3][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[3][9] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[3][9] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[3][9] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[3][9] .mask = 16'hCC00;
defparam \macro_inst|controller|sm_pwm|pwmList[3][9] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[3][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[3][9] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[40][0]~75_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][0] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[40][0] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][0] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[40][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[40][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[40][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan81~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(SyncReset_X60_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan81~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][10] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[40][10] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][10] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[40][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[40][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[40][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan81~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(SyncReset_X60_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan81~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][11] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[40][11] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][11] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[40][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[40][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[40][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan81~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(SyncReset_X60_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan81~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][12] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[40][12] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][12] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[40][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[40][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[40][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan81~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(SyncReset_X60_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan81~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][13] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[40][13] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][13] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[40][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[40][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[40][14]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan81~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(SyncReset_X60_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y10_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan81~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][14] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[40][14] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][14] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[40][14] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[40][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][15] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[40][7]~q ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X62_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ),
	.SyncReset(SyncReset_X62_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y9_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~242_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][15] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[40][15] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][15] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[40][15] .mask = 16'hFF72;
defparam \macro_inst|controller|sm_pwm|pwmList[40][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[40][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan82~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X62_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ),
	.SyncReset(SyncReset_X62_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan82~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][1] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[40][1] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][1] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[40][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[40][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[40][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan82~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X62_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ),
	.SyncReset(SyncReset_X62_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan82~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][2] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[40][2] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][2] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[40][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[40][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[40][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan82~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X62_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ),
	.SyncReset(SyncReset_X62_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan82~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][3] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[40][3] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][3] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[40][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[40][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[40][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan82~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X62_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ),
	.SyncReset(SyncReset_X62_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan82~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][4] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[40][4] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][4] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[40][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[40][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X62_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[40][5]~74_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][5] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[40][5] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][5] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[40][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[40][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan82~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X62_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y9_SIG ),
	.SyncReset(SyncReset_X62_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y9_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan82~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][6] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[40][6] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][6] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[40][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[40][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[40][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][7] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[40][7] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][7] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[40][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[40][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[40][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(SyncReset_X60_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan81~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][8] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[40][8] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][8] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[40][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[40][9] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[40][9]~q ),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan81~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[40][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~66_combout_X60_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y10_SIG ),
	.SyncReset(SyncReset_X60_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan81~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[40][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[40][9] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[40][9] .coord_y = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[40][9] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][9] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[40][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[40][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[40][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X60_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[41][0]~27_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][0] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[41][0] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[41][0] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[41][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[41][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[41][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan83~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X61_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y10_SIG ),
	.SyncReset(SyncReset_X61_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan83~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][10] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[41][10] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[41][10] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[41][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[41][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][11] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[41][11]~q ),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan83~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X61_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y10_SIG ),
	.SyncReset(SyncReset_X61_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan83~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][11] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[41][11] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[41][11] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[41][11] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[41][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[41][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan83~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X61_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y10_SIG ),
	.SyncReset(SyncReset_X61_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan83~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][12] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[41][12] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[41][12] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[41][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[41][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[41][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan83~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X61_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y10_SIG ),
	.SyncReset(SyncReset_X61_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan83~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][13] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[41][13] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[41][13] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[41][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[41][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][14] (
	.A(\macro_inst|controller|sm_pwm|pwmList[41][0]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X60_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ),
	.SyncReset(SyncReset_X60_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan84~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][14] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[41][14] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[41][14] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[41][14] .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|pwmList[41][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][14] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[10][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan21~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X61_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y10_SIG ),
	.SyncReset(SyncReset_X61_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan21~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][15] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[41][15] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[41][15] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[41][15] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[41][15] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][15] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[41][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan84~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X60_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ),
	.SyncReset(SyncReset_X60_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan84~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][1] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[41][1] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[41][1] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[41][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[41][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[41][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan84~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X60_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ),
	.SyncReset(SyncReset_X60_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan84~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][2] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[41][2] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[41][2] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[41][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[41][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[41][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan84~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X60_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ),
	.SyncReset(SyncReset_X60_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan84~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][3] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[41][3] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[41][3] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[41][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[41][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[41][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan84~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X60_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ),
	.SyncReset(SyncReset_X60_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan84~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][4] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[41][4] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[41][4] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[41][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[41][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][5] (
	.A(vcc),
	.B(\rv32.mem_ahb_hwdata[5] ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X60_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[41][5]~26_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][5] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[41][5] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[41][5] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[41][5] .mask = 16'h3333;
defparam \macro_inst|controller|sm_pwm|pwmList[41][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][6] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[41][6]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan84~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X60_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ),
	.SyncReset(SyncReset_X60_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y6_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan84~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][6] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[41][6] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[41][6] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[41][6] .mask = 16'h5F05;
defparam \macro_inst|controller|sm_pwm|pwmList[41][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][7] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[41][5]~q ),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan84~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X60_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y6_SIG ),
	.SyncReset(SyncReset_X60_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan84~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][7] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[41][7] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[41][7] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[41][7] .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|pwmList[41][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][7] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][8] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[41][8]~q ),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X61_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y10_SIG ),
	.SyncReset(SyncReset_X61_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan83~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][8] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[41][8] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[41][8] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][8] .mask = 16'h0044;
defparam \macro_inst|controller|sm_pwm|pwmList[41][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[41][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[41][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan83~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[41][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~36_combout_X61_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y10_SIG ),
	.SyncReset(SyncReset_X61_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan83~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[41][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[41][9] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[41][9] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[41][9] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[41][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[41][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[41][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[42][0]~77_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][0] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[42][0] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[42][0] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[42][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[42][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[42][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan85~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(SyncReset_X62_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan85~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][10] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[42][10] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[42][10] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[42][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[42][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[42][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan85~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(SyncReset_X62_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan85~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][11] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[42][11] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[42][11] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[42][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[42][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[42][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan85~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(SyncReset_X62_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan85~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][12] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[42][12] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[42][12] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[42][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[42][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[42][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan85~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(SyncReset_X62_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan85~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][13] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[42][13] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[42][13] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[42][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[42][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][14] (
	.A(\macro_inst|controller|sm_pwm|pwmList[42][14]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan85~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(SyncReset_X62_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y11_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan85~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][14] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[42][14] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[42][14] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[42][14] .mask = 16'h2B2B;
defparam \macro_inst|controller|sm_pwm|pwmList[42][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][15] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[42][7]~q ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|LessThan86~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ),
	.SyncReset(SyncReset_X62_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~244_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][15] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[42][15] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[42][15] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[42][15] .mask = 16'h72FA;
defparam \macro_inst|controller|sm_pwm|pwmList[42][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][1] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[42][1]~q ),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan86~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ),
	.SyncReset(SyncReset_X62_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan86~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][1] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[42][1] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[42][1] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[42][1] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[42][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[42][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan86~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ),
	.SyncReset(SyncReset_X62_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan86~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][2] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[42][2] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[42][2] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[42][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[42][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][3] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[42][3]~q ),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan86~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ),
	.SyncReset(SyncReset_X62_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan86~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][3] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[42][3] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[42][3] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[42][3] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[42][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[42][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan86~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ),
	.SyncReset(SyncReset_X62_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y7_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan86~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][4] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[42][4] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[42][4] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[42][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[42][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[42][5]~76_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][5] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[42][5] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[42][5] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[42][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[42][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan86~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ),
	.SyncReset(SyncReset_X62_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan86~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][6] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[42][6] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[42][6] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[42][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[42][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][7] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|LessThan85~12_combout ),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[42][15]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y7_SIG ),
	.SyncReset(SyncReset_X62_Y7_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y7_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~196_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][7] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[42][7] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[42][7] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[42][7] .mask = 16'hAF27;
defparam \macro_inst|controller|sm_pwm|pwmList[42][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[42][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(SyncReset_X62_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan85~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][8] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[42][8] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[42][8] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[42][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[42][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[42][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[42][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan85~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[42][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~68_combout_X62_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y11_SIG ),
	.SyncReset(SyncReset_X62_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X62_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan85~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[42][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[42][9] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[42][9] .coord_y = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[42][9] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[42][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[42][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[42][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[42][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X59_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[43][0]~29_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][0] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[43][0] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[43][0] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[43][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[43][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[43][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan87~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X60_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ),
	.SyncReset(SyncReset_X60_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan87~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][10] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[43][10] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[43][10] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[43][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[43][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[43][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan87~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X60_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ),
	.SyncReset(SyncReset_X60_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan87~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][11] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[43][11] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[43][11] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[43][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[43][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][12] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[43][12]~q ),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan87~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X60_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ),
	.SyncReset(SyncReset_X60_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan87~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][12] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[43][12] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[43][12] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[43][12] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[43][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[43][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan87~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X60_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ),
	.SyncReset(SyncReset_X60_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan87~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][13] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[43][13] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[43][13] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[43][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[43][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[43][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan87~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X60_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ),
	.SyncReset(SyncReset_X60_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y12_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan87~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][14] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[43][14] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[43][14] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[43][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[43][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][15] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[15] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X59_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[43][15]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][15] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[43][15] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[43][15] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[43][15] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[43][15] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][15] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[43][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan88~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X59_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ),
	.SyncReset(SyncReset_X59_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan88~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][1] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[43][1] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[43][1] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[43][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[43][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[43][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan88~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X59_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ),
	.SyncReset(SyncReset_X59_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan88~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][2] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[43][2] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[43][2] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[43][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[43][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[43][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan88~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X59_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ),
	.SyncReset(SyncReset_X59_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan88~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][3] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[43][3] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[43][3] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[43][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[43][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[43][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan88~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X59_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ),
	.SyncReset(SyncReset_X59_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan88~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][4] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[43][4] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[43][4] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[43][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[43][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X59_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[43][5]~28_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][5] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[43][5] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[43][5] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[43][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[43][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan88~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X59_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ),
	.SyncReset(SyncReset_X59_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y10_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan88~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][6] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[43][6] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[43][6] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[43][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[43][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][7] (
	.A(\macro_inst|controller|sm_pwm|pwmList[43][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan88~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X59_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y10_SIG ),
	.SyncReset(SyncReset_X59_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan88~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][7] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[43][7] .coord_y = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[43][7] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[43][7] .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|pwmList[43][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][7] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[43][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X60_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ),
	.SyncReset(SyncReset_X60_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan87~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][8] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[43][8] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[43][8] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[43][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[43][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[43][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[43][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan87~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[43][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~38_combout_X60_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y12_SIG ),
	.SyncReset(SyncReset_X60_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan87~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[43][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[43][9] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[43][9] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[43][9] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[43][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[43][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[43][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[43][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][0] (
	.A(\rv32.mem_ahb_hwdata[0] ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X59_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[44][0]~79_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][0] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[44][0] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][0] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[44][0] .mask = 16'h5555;
defparam \macro_inst|controller|sm_pwm|pwmList[44][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[44][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan89~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan89~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][10] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[44][10] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][10] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[44][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[44][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[44][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan89~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan89~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][11] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[44][11] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][11] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[44][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[44][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[44][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan89~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan89~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][12] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[44][12] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][12] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[44][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[44][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[44][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan89~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan89~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][13] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[44][13] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][13] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[44][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[44][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[44][14]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan89~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan89~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][14] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[44][14] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][14] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[44][14] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[44][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[44][7]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|LessThan90~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X59_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ),
	.SyncReset(SyncReset_X59_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y5_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~246_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][15] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[44][15] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][15] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[44][15] .mask = 16'h74FC;
defparam \macro_inst|controller|sm_pwm|pwmList[44][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[44][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan90~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X59_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ),
	.SyncReset(SyncReset_X59_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan90~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][1] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[44][1] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][1] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[44][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[44][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[44][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan90~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X59_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ),
	.SyncReset(SyncReset_X59_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan90~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][2] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[44][2] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][2] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[44][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[44][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][3] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X59_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ),
	.SyncReset(SyncReset_X59_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y5_VCC),
	.LutOut(\macro_inst|mem_ahb_hrdata[3]~3_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][3] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[44][3] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][3] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[44][3] .mask = 16'hCC00;
defparam \macro_inst|controller|sm_pwm|pwmList[44][3] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][3] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[44][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan90~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X59_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ),
	.SyncReset(SyncReset_X59_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y5_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan90~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][4] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[44][4] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][4] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[44][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[44][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][5] (
	.A(vcc),
	.B(\rv32.mem_ahb_hwdata[5] ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X59_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[44][5]~78_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][5] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[44][5] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][5] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[44][5] .mask = 16'h3333;
defparam \macro_inst|controller|sm_pwm|pwmList[44][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[44][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan90~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X59_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ),
	.SyncReset(SyncReset_X59_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y5_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan90~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][6] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[44][6] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][6] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[44][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[44][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][7] (
	.A(\macro_inst|controller|sm_pwm|pwmList[44][15]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|LessThan89~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X59_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y5_SIG ),
	.SyncReset(SyncReset_X59_Y5_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y5_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~198_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][7] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[44][7] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][7] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[44][7] .mask = 16'h8BCF;
defparam \macro_inst|controller|sm_pwm|pwmList[44][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[44][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan89~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][8] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[44][8] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][8] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[44][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[44][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[44][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan89~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[44][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~69_combout_X60_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y4_SIG ),
	.SyncReset(SyncReset_X60_Y4_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y4_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan89~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[44][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[44][9] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[44][9] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[44][9] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[44][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[44][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[44][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X58_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[45][0]~31_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][0] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[45][0] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[45][0] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[45][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[45][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan91~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X57_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y6_SIG ),
	.SyncReset(SyncReset_X57_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan91~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][10] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[45][10] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[45][10] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[45][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[45][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][11] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[45][11]~q ),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan91~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X57_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y6_SIG ),
	.SyncReset(SyncReset_X57_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan91~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][11] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[45][11] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[45][11] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[45][11] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[45][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[45][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan91~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X57_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y6_SIG ),
	.SyncReset(SyncReset_X57_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan91~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][12] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[45][12] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[45][12] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[45][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[45][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[45][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan91~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X57_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y6_SIG ),
	.SyncReset(SyncReset_X57_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan91~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][13] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[45][13] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[45][13] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[45][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[45][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][14] (
	.A(\macro_inst|controller|sm_pwm|pwmList[45][14]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan91~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X57_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y6_SIG ),
	.SyncReset(SyncReset_X57_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y6_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan91~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][14] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[45][14] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[45][14] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[45][14] .mask = 16'h2B2B;
defparam \macro_inst|controller|sm_pwm|pwmList[45][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][15] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[15] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X57_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[45][15]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][15] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[45][15] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[45][15] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][15] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[45][15] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][15] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][1] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[45][1]~q ),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan92~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X58_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y10_SIG ),
	.SyncReset(SyncReset_X58_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan92~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][1] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[45][1] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[45][1] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[45][1] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[45][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[45][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan92~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X58_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y10_SIG ),
	.SyncReset(SyncReset_X58_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan92~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][2] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[45][2] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[45][2] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[45][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[45][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[45][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan92~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X58_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y10_SIG ),
	.SyncReset(SyncReset_X58_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan92~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][3] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[45][3] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[45][3] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[45][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[45][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[45][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan92~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X58_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y10_SIG ),
	.SyncReset(SyncReset_X58_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan92~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][4] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[45][4] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[45][4] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[45][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[45][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X57_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[45][5]~30_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][5] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[45][5] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[45][5] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[45][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[45][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[45][6]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan92~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X58_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y10_SIG ),
	.SyncReset(SyncReset_X58_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y10_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan92~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][6] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[45][6] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[45][6] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[45][6] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[45][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X57_Y7_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y7_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[45][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][7] .coord_x = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[45][7] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[45][7] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[45][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[45][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[45][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X57_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y6_SIG ),
	.SyncReset(SyncReset_X57_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan91~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][8] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[45][8] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[45][8] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[45][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[45][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[45][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[45][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan91~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[45][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~39_combout_X57_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y6_SIG ),
	.SyncReset(SyncReset_X57_Y6_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y6_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan91~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[45][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[45][9] .coord_x = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[45][9] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[45][9] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[45][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[45][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[45][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[45][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[46][0]~81_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][0] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[46][0] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][0] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[46][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[46][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[46][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan93~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(SyncReset_X58_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan93~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][10] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[46][10] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][10] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[46][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[46][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[46][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan93~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(SyncReset_X58_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan93~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][11] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[46][11] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][11] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[46][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[46][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[46][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan93~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(SyncReset_X58_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan93~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][12] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[46][12] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][12] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[46][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[46][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[46][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan93~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(SyncReset_X58_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan93~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][13] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[46][13] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][13] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[46][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[46][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[46][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan93~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(SyncReset_X58_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y1_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan93~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][14] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[46][14] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][14] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[46][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[46][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][15] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[15] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X57_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[46][15]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][15] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[46][15] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[46][15] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[46][15] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[46][15] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][15] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][1] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[46][1]~q ),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan94~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X57_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y1_SIG ),
	.SyncReset(SyncReset_X57_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan94~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][1] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[46][1] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[46][1] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[46][1] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[46][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][2] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.B(\macro_inst|controller|sm_pwm|pwmList[46][2]~q ),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan94~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X57_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y1_SIG ),
	.SyncReset(SyncReset_X57_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan94~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][2] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[46][2] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[46][2] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[46][2] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[46][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[46][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan94~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X57_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y1_SIG ),
	.SyncReset(SyncReset_X57_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan94~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][3] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[46][3] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[46][3] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[46][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[46][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[46][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan94~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X57_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y1_SIG ),
	.SyncReset(SyncReset_X57_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan94~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][4] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[46][4] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[46][4] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[46][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[46][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X57_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[46][5]~80_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][5] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[46][5] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[46][5] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[46][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[46][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan94~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X57_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y1_SIG ),
	.SyncReset(SyncReset_X57_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y1_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan94~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][6] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[46][6] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[46][6] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[46][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[46][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X57_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[46][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][7] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[46][7] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[46][7] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[46][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[46][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[46][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(SyncReset_X58_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan93~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][8] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[46][8] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][8] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[46][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[46][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[46][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan93~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[46][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~70_combout_X58_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y1_SIG ),
	.SyncReset(SyncReset_X58_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan93~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[46][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[46][9] .coord_x = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[46][9] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][9] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[46][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[46][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[46][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X60_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[47][0]~33_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][0] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[47][0] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][0] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[47][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[47][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][10] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[47][0]~q ),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X60_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(SyncReset_X60_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan96~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][10] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[47][10] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][10] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[47][10] .mask = 16'h0011;
defparam \macro_inst|controller|sm_pwm|pwmList[47][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[47][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan95~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X61_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ),
	.SyncReset(SyncReset_X61_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan95~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][11] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[47][11] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][11] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[47][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[47][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[47][5]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan96~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X60_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(SyncReset_X60_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan96~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][12] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[47][12] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][12] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[47][12] .mask = 16'h008E;
defparam \macro_inst|controller|sm_pwm|pwmList[47][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[47][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan95~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X61_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ),
	.SyncReset(SyncReset_X61_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan95~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][13] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[47][13] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][13] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[47][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[47][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[47][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan95~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X61_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ),
	.SyncReset(SyncReset_X61_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y1_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan95~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][14] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[47][14] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][14] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[47][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[47][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[47][7]~q ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|LessThan96~12_combout ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X60_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(SyncReset_X60_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y1_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~104_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][15] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[47][15] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][15] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[47][15] .mask = 16'h74FC;
defparam \macro_inst|controller|sm_pwm|pwmList[47][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[47][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan96~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X60_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(SyncReset_X60_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan96~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][1] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[47][1] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][1] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[47][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[47][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[47][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan96~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X60_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(SyncReset_X60_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan96~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][2] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[47][2] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][2] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[47][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[47][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[47][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan96~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X60_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(SyncReset_X60_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan96~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][3] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[47][3] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][3] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[47][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[47][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[47][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan96~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X60_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(SyncReset_X60_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan96~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][4] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[47][4] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][4] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[47][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[47][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X60_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[47][5]~32_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][5] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[47][5] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][5] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[47][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[47][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan96~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X60_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(SyncReset_X60_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y1_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan96~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][6] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[47][6] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][6] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[47][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[47][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][7] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|LessThan95~12_combout ),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[47][15]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X60_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y1_SIG ),
	.SyncReset(SyncReset_X60_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y1_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~56_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][7] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[47][7] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][7] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[47][7] .mask = 16'hAF27;
defparam \macro_inst|controller|sm_pwm|pwmList[47][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][8] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[47][8]~q ),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X61_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ),
	.SyncReset(SyncReset_X61_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan95~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][8] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[47][8] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][8] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[47][8] .mask = 16'h0044;
defparam \macro_inst|controller|sm_pwm|pwmList[47][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[47][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[47][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan95~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[47][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~40_combout_X61_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y1_SIG ),
	.SyncReset(SyncReset_X61_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan95~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[47][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[47][9] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[47][9] .coord_y = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][9] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[47][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[47][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[47][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[47][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[4][0]~73_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][0] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[4][0] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[4][0] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[4][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[4][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[4][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan9~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(SyncReset_X57_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan9~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][10] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[4][10] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[4][10] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[4][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[4][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][11] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[4][11]~q ),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan9~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(SyncReset_X57_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan9~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][11] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[4][11] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[4][11] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[4][11] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[4][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[4][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan9~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(SyncReset_X57_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan9~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][12] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[4][12] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[4][12] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[4][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[4][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[4][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan9~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(SyncReset_X57_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan9~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][13] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[4][13] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[4][13] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[4][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[4][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][14] (
	.A(\macro_inst|controller|sm_pwm|pwmList[4][14]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan9~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(SyncReset_X57_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y10_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan9~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][14] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[4][14] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[4][14] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[4][14] .mask = 16'h2B2B;
defparam \macro_inst|controller|sm_pwm|pwmList[4][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][15] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|LessThan10~12_combout ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[4][7]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y12_SIG ),
	.SyncReset(SyncReset_X57_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y12_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~240_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][15] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[4][15] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[4][15] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[4][15] .mask = 16'h72FA;
defparam \macro_inst|controller|sm_pwm|pwmList[4][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[4][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan10~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y12_SIG ),
	.SyncReset(SyncReset_X57_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan10~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][1] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[4][1] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[4][1] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[4][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[4][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[4][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan10~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y12_SIG ),
	.SyncReset(SyncReset_X57_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan10~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][2] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[4][2] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[4][2] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[4][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[4][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[4][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan10~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y12_SIG ),
	.SyncReset(SyncReset_X57_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan10~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][3] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[4][3] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[4][3] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[4][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[4][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[4][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan10~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y12_SIG ),
	.SyncReset(SyncReset_X57_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan10~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][4] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[4][4] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[4][4] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[4][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[4][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X58_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[4][5]~72_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][5] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[4][5] .coord_y = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[4][5] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[4][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[4][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[4][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan10~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y12_SIG ),
	.SyncReset(SyncReset_X57_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y12_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan10~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][6] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[4][6] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[4][6] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[4][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[4][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y12_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[4][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][7] .coord_x = 18;
defparam \macro_inst|controller|sm_pwm|pwmList[4][7] .coord_y = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[4][7] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[4][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[4][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[4][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(SyncReset_X57_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan9~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][8] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[4][8] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[4][8] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[4][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[4][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[4][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan9~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[4][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~65_combout_X57_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y10_SIG ),
	.SyncReset(SyncReset_X57_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan9~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[4][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[4][9] .coord_x = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[4][9] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[4][9] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[4][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[4][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[4][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X59_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[5][0]~25_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][0] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][0] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[5][0] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[5][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[5][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[5][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan11~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X60_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ),
	.SyncReset(SyncReset_X60_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan11~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][10] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][10] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[5][10] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[5][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[5][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][11] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[5][11]~q ),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan11~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X60_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ),
	.SyncReset(SyncReset_X60_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan11~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][11] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][11] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[5][11] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[5][11] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[5][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[5][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan11~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X60_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ),
	.SyncReset(SyncReset_X60_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan11~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][12] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][12] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[5][12] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[5][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[5][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][13] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[5][13]~q ),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan11~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X60_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ),
	.SyncReset(SyncReset_X60_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan11~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][13] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][13] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[5][13] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[5][13] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[5][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[5][14]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan11~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X60_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ),
	.SyncReset(SyncReset_X60_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y11_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan11~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][14] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][14] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[5][14] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[5][14] .mask = 16'h3F03;
defparam \macro_inst|controller|sm_pwm|pwmList[5][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][15] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[15] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X59_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[5][15]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][15] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][15] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[5][15] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][15] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[5][15] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][15] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[5][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan12~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X59_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y11_SIG ),
	.SyncReset(SyncReset_X59_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan12~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][1] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][1] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[5][1] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[5][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[5][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[5][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan12~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X59_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y11_SIG ),
	.SyncReset(SyncReset_X59_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan12~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][2] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][2] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[5][2] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[5][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[5][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][3] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[5][3]~q ),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan12~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X59_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y11_SIG ),
	.SyncReset(SyncReset_X59_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan12~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][3] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][3] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[5][3] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[5][3] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[5][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[5][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan12~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X59_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y11_SIG ),
	.SyncReset(SyncReset_X59_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan12~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][4] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][4] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[5][4] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[5][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[5][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X59_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[5][5]~24_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][5] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][5] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[5][5] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[5][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[5][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[5][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan12~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X59_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y11_SIG ),
	.SyncReset(SyncReset_X59_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y11_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan12~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][6] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][6] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[5][6] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[5][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[5][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X59_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[5][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][7] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][7] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[5][7] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[5][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[5][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][8] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[5][8]~q ),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X60_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ),
	.SyncReset(SyncReset_X60_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan11~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][8] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][8] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[5][8] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[5][8] .mask = 16'h0044;
defparam \macro_inst|controller|sm_pwm|pwmList[5][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[5][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[5][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan11~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[5][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~34_combout_X60_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ),
	.SyncReset(SyncReset_X60_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan11~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[5][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[5][9] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[5][9] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[5][9] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[5][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[5][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[5][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[5][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X59_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[6][0]~83_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][0] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][0] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[6][0] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[6][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[6][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[6][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan13~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X58_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ),
	.SyncReset(SyncReset_X58_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan13~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][10] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][10] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[6][10] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[6][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[6][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[6][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan13~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X58_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ),
	.SyncReset(SyncReset_X58_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan13~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][11] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][11] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[6][11] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[6][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[6][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[6][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan13~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X58_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ),
	.SyncReset(SyncReset_X58_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan13~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][12] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][12] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[6][12] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[6][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[6][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][13] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[6][13]~q ),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan13~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X58_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ),
	.SyncReset(SyncReset_X58_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan13~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][13] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][13] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[6][13] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[6][13] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[6][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[6][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan13~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X58_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ),
	.SyncReset(SyncReset_X58_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y2_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan13~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][14] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][14] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[6][14] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[6][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[6][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][15] (
	.A(\macro_inst|controller|sm_pwm|pwmList[6][7]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X59_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ),
	.SyncReset(SyncReset_X59_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y1_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~250_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][15] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][15] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[6][15] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[6][15] .mask = 16'hDDFC;
defparam \macro_inst|controller|sm_pwm|pwmList[6][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[6][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan14~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X59_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ),
	.SyncReset(SyncReset_X59_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan14~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][1] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][1] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[6][1] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[6][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[6][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][2] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.B(\macro_inst|controller|sm_pwm|pwmList[6][2]~q ),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan14~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X59_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ),
	.SyncReset(SyncReset_X59_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan14~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][2] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][2] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[6][2] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[6][2] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[6][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[6][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan14~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X59_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ),
	.SyncReset(SyncReset_X59_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan14~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][3] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][3] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[6][3] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[6][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[6][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[6][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan14~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X59_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ),
	.SyncReset(SyncReset_X59_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y1_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan14~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][4] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][4] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[6][4] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[6][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[6][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X59_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[6][5]~82_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][5] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][5] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[6][5] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[6][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[6][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[6][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan14~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X59_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ),
	.SyncReset(SyncReset_X59_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y1_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan14~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][6] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][6] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[6][6] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[6][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[6][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][7] (
	.A(\macro_inst|controller|sm_pwm|LessThan13~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[6][15]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X59_Y1_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y1_SIG ),
	.SyncReset(SyncReset_X59_Y1_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X59_Y1_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~202_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][7] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][7] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[6][7] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][7] .mask = 16'hCF47;
defparam \macro_inst|controller|sm_pwm|pwmList[6][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[6][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X58_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ),
	.SyncReset(SyncReset_X58_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan13~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][8] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][8] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[6][8] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[6][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[6][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[6][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan13~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[6][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~72_combout_X58_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y2_SIG ),
	.SyncReset(SyncReset_X58_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y2_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan13~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[6][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[6][9] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[6][9] .coord_y = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[6][9] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[6][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[6][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[6][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X62_Y6_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X62_Y6_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[7][0]~35_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][0] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[7][0] .coord_y = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[7][0] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[7][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[7][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[7][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan15~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan15~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][10] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[7][10] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][10] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[7][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[7][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[7][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan15~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan15~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][11] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[7][11] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][11] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[7][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[7][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[7][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan15~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan15~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][12] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[7][12] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][12] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[7][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[7][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][13] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[7][13]~q ),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan15~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan15~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][13] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[7][13] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][13] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[7][13] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[7][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[7][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan15~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan15~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][14] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[7][14] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][14] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[7][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][15] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[15] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[7][15]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][15] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[7][15] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][15] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][15] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[7][15] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][15] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[7][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan16~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X58_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y10_SIG ),
	.SyncReset(SyncReset_X58_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan16~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][1] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[7][1] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][1] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[7][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[7][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[7][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan16~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X58_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y10_SIG ),
	.SyncReset(SyncReset_X58_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan16~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][2] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[7][2] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][2] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[7][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[7][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[7][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan16~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X58_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y10_SIG ),
	.SyncReset(SyncReset_X58_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan16~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][3] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[7][3] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][3] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[7][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[7][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][4] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.B(\macro_inst|controller|sm_pwm|pwmList[7][4]~q ),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan16~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X58_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y10_SIG ),
	.SyncReset(SyncReset_X58_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y10_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan16~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][4] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[7][4] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][4] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[7][4] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[7][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X58_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y10_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[7][5]~34_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][5] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[7][5] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][5] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[7][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[7][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[7][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan16~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X58_Y10_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y10_SIG ),
	.SyncReset(SyncReset_X58_Y10_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y10_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan16~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][6] .coord_x = 17;
defparam \macro_inst|controller|sm_pwm|pwmList[7][6] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][6] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[7][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][7] (
	.A(\macro_inst|controller|sm_pwm|pwmList[7][15]~q ),
	.B(\macro_inst|controller|sm_pwm|LessThan15~12_combout ),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~58_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][7] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[7][7] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][7] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[7][7] .mask = 16'hBB0F;
defparam \macro_inst|controller|sm_pwm|pwmList[7][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[7][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan15~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][8] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[7][8] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][8] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[7][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[7][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[7][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan15~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[7][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~42_combout_X60_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y8_SIG ),
	.SyncReset(SyncReset_X60_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan15~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[7][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[7][9] .coord_x = 16;
defparam \macro_inst|controller|sm_pwm|pwmList[7][9] .coord_y = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[7][9] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[7][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[7][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[7][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[7][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X61_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[8][0]~85_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][0] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][0] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[8][0] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[8][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[8][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[8][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan17~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X60_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ),
	.SyncReset(SyncReset_X60_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan17~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][10] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][10] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[8][10] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[8][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[8][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][11] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.B(\macro_inst|controller|sm_pwm|pwmList[8][11]~q ),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan17~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X60_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ),
	.SyncReset(SyncReset_X60_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan17~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][11] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][11] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[8][11] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[8][11] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[8][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[8][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan17~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X60_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ),
	.SyncReset(SyncReset_X60_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan17~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][12] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][12] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[8][12] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[8][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[8][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][13] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.B(\macro_inst|controller|sm_pwm|pwmList[8][13]~q ),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan17~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X60_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ),
	.SyncReset(SyncReset_X60_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan17~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][13] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][13] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[8][13] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[8][13] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[8][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[8][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan17~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X60_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ),
	.SyncReset(SyncReset_X60_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y11_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan17~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][14] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][14] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[8][14] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[8][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[8][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][15] (
	.A(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[8][7]~q ),
	.C(\rv32.mem_ahb_hwdata[15] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [7]),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X61_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ),
	.SyncReset(SyncReset_X61_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y8_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~204_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][15] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][15] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[8][15] .coord_z = 15;
defparam \macro_inst|controller|sm_pwm|pwmList[8][15] .mask = 16'hFFB1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][15] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][15] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][15] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][1] (
	.A(\macro_inst|controller|sm_pwm|pwmList[8][1]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan18~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X61_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ),
	.SyncReset(SyncReset_X61_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan18~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][1] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][1] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[8][1] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[8][1] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[8][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[8][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan18~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X61_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ),
	.SyncReset(SyncReset_X61_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan18~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][2] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][2] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[8][2] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[8][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[8][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[8][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan18~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X61_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ),
	.SyncReset(SyncReset_X61_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan18~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][3] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][3] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[8][3] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[8][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[8][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[8][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan18~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X61_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ),
	.SyncReset(SyncReset_X61_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y8_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan18~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][4] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][4] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[8][4] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[8][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[8][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][5] (
	.A(vcc),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[5] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X61_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[8][5]~84_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][5] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][5] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[8][5] .coord_z = 14;
defparam \macro_inst|controller|sm_pwm|pwmList[8][5] .mask = 16'h0F0F;
defparam \macro_inst|controller|sm_pwm|pwmList[8][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][6] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.B(vcc),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[8][6]~q ),
	.Cin(\macro_inst|controller|sm_pwm|LessThan18~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X61_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ),
	.SyncReset(SyncReset_X61_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y8_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan18~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][6] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][6] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[8][6] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[8][6] .mask = 16'h5F05;
defparam \macro_inst|controller|sm_pwm|pwmList[8][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][7] (
	.A(\macro_inst|controller|sm_pwm|LessThan18~12_combout ),
	.B(\macro_inst|controller|sm_pwm|motor_flags [0]),
	.C(\rv32.mem_ahb_hwdata[7] ),
	.D(\macro_inst|controller|sm_pwm|pwmList[8][15]~q ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X61_Y8_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X61_Y8_SIG ),
	.SyncReset(SyncReset_X61_Y8_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X61_Y8_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|data~252_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][7] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][7] .coord_y = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[8][7] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][7] .mask = 16'h7F4C;
defparam \macro_inst|controller|sm_pwm|pwmList[8][7] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][7] .FeedbackMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][7] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][8] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.B(\macro_inst|controller|sm_pwm|pwmList[8][8]~q ),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X60_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ),
	.SyncReset(SyncReset_X60_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan17~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][8] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][8] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[8][8] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[8][8] .mask = 16'h0044;
defparam \macro_inst|controller|sm_pwm|pwmList[8][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[8][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[8][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan17~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[8][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~73_combout_X60_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y11_SIG ),
	.SyncReset(SyncReset_X60_Y11_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y11_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan17~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[8][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[8][9] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[8][9] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[8][9] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[8][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[8][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[8][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[8][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[0] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[9][0]~37_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][0]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][0] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[9][0] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[9][0] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][0] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[9][0] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][0] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][0] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][0] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][10] (
	.A(\macro_inst|controller|sm_pwm|pwmList[9][10]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[10] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan19~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][10]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(SyncReset_X60_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan19~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][10]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][10] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[9][10] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[9][10] .coord_z = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[9][10] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[9][10] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][10] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][10] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][10] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][10] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][11] (
	.A(\macro_inst|controller|sm_pwm|pwmList[9][11]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[11] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan19~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][11]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(SyncReset_X60_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan19~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][11]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][11] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[9][11] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[9][11] .coord_z = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[9][11] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[9][11] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][11] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][11] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][11] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][11] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][12] (
	.A(\macro_inst|controller|sm_pwm|pwmList[9][12]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[12] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan19~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][12]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(SyncReset_X60_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan19~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][12]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][12] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[9][12] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[9][12] .coord_z = 5;
defparam \macro_inst|controller|sm_pwm|pwmList[9][12] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[9][12] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][12] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][12] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][12] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][12] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][13] (
	.A(\macro_inst|controller|sm_pwm|pwmList[9][13]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [5]),
	.C(\rv32.mem_ahb_hwdata[13] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan19~9_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][13]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(SyncReset_X60_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan19~11_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][13]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][13] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[9][13] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[9][13] .coord_z = 6;
defparam \macro_inst|controller|sm_pwm|pwmList[9][13] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[9][13] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][13] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][13] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][13] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][13] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][14] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[9][14]~q ),
	.C(\rv32.mem_ahb_hwdata[14] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan19~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][14]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(SyncReset_X60_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y9_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan19~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][14]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][14] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[9][14] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[9][14] .coord_z = 7;
defparam \macro_inst|controller|sm_pwm|pwmList[9][14] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[9][14] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][14] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][14] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][14] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][14] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][15] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[15] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][15]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X59_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[9][15]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][15]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][15] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[9][15] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[9][15] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[9][15] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[9][15] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][15] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][15] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][15] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][15] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][1] (
	.A(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.B(\macro_inst|controller|sm_pwm|pwmList[9][1]~q ),
	.C(\rv32.mem_ahb_hwdata[1] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan20~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X58_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y12_SIG ),
	.SyncReset(SyncReset_X58_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan20~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][1]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][1] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[9][1] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[9][1] .coord_z = 8;
defparam \macro_inst|controller|sm_pwm|pwmList[9][1] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[9][1] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][1] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][1] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][1] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][1] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][2] (
	.A(\macro_inst|controller|sm_pwm|pwmList[9][2]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [2]),
	.C(\rv32.mem_ahb_hwdata[2] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan20~3_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X58_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y12_SIG ),
	.SyncReset(SyncReset_X58_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan20~5_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][2]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][2] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[9][2] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[9][2] .coord_z = 9;
defparam \macro_inst|controller|sm_pwm|pwmList[9][2] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[9][2] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][2] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][2] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][2] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][2] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][3] (
	.A(\macro_inst|controller|sm_pwm|pwmList[9][3]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [3]),
	.C(\rv32.mem_ahb_hwdata[3] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan20~5_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X58_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y12_SIG ),
	.SyncReset(SyncReset_X58_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan20~7_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][3]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][3] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[9][3] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[9][3] .coord_z = 10;
defparam \macro_inst|controller|sm_pwm|pwmList[9][3] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[9][3] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][3] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][3] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][3] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][3] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][4] (
	.A(\macro_inst|controller|sm_pwm|pwmList[9][4]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [4]),
	.C(\rv32.mem_ahb_hwdata[4] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan20~7_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X58_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y12_SIG ),
	.SyncReset(SyncReset_X58_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y12_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan20~9_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][4]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][4] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[9][4] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[9][4] .coord_z = 11;
defparam \macro_inst|controller|sm_pwm|pwmList[9][4] .mask = 16'h002B;
defparam \macro_inst|controller|sm_pwm|pwmList[9][4] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][4] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][4] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][4] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][4] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[5] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X59_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[9][5]~36_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][5]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][5] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[9][5] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[9][5] .coord_z = 0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][5] .mask = 16'h00FF;
defparam \macro_inst|controller|sm_pwm|pwmList[9][5] .modeMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][5] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][5] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][5] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][6] (
	.A(vcc),
	.B(\macro_inst|controller|sm_pwm|pwmList[9][6]~q ),
	.C(\rv32.mem_ahb_hwdata[6] ),
	.D(\macro_inst|controller|sm_pwm|pwmCnt [6]),
	.Cin(\macro_inst|controller|sm_pwm|LessThan20~11_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X58_Y12_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X58_Y12_SIG ),
	.SyncReset(SyncReset_X58_Y12_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X58_Y12_VCC),
	.LutOut(\macro_inst|controller|sm_pwm|LessThan20~12_combout ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][6]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][6] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[9][6] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[9][6] .coord_z = 13;
defparam \macro_inst|controller|sm_pwm|pwmList[9][6] .mask = 16'h0CCF;
defparam \macro_inst|controller|sm_pwm|pwmList[9][6] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][6] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][6] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][6] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][7] (
	.A(),
	.B(),
	.C(vcc),
	.D(\rv32.mem_ahb_hwdata[7] ),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X59_Y11_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X59_Y11_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|controller|sm_pwm|pwmList[9][7]__feeder__LutOut ),
	.Cout(),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][7]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][7] .coord_x = 19;
defparam \macro_inst|controller|sm_pwm|pwmList[9][7] .coord_y = 3;
defparam \macro_inst|controller|sm_pwm|pwmList[9][7] .coord_z = 12;
defparam \macro_inst|controller|sm_pwm|pwmList[9][7] .mask = 16'hFF00;
defparam \macro_inst|controller|sm_pwm|pwmList[9][7] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][7] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][7] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][7] .BypassEn = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][8] (
	.A(\macro_inst|controller|sm_pwm|pwmList[9][8]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [0]),
	.C(\rv32.mem_ahb_hwdata[8] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][8]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(SyncReset_X60_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan19~1_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][8]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][8] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[9][8] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[9][8] .coord_z = 1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][8] .mask = 16'h0022;
defparam \macro_inst|controller|sm_pwm|pwmList[9][8] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][8] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][8] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][8] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][8] .CarryEnb = 1'b0;

alta_slice \macro_inst|controller|sm_pwm|pwmList[9][9] (
	.A(\macro_inst|controller|sm_pwm|pwmList[9][9]~q ),
	.B(\macro_inst|controller|sm_pwm|pwmCnt [1]),
	.C(\rv32.mem_ahb_hwdata[9] ),
	.D(vcc),
	.Cin(\macro_inst|controller|sm_pwm|LessThan19~1_cout ),
	.Qin(\macro_inst|controller|sm_pwm|pwmList[9][9]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|controller|sm_pwm|Decoder0~43_combout_X60_Y9_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X60_Y9_SIG ),
	.SyncReset(SyncReset_X60_Y9_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X60_Y9_VCC),
	.LutOut(),
	.Cout(\macro_inst|controller|sm_pwm|LessThan19~3_cout ),
	.Q(\macro_inst|controller|sm_pwm|pwmList[9][9]~q ));
defparam \macro_inst|controller|sm_pwm|pwmList[9][9] .coord_x = 20;
defparam \macro_inst|controller|sm_pwm|pwmList[9][9] .coord_y = 4;
defparam \macro_inst|controller|sm_pwm|pwmList[9][9] .coord_z = 2;
defparam \macro_inst|controller|sm_pwm|pwmList[9][9] .mask = 16'h004D;
defparam \macro_inst|controller|sm_pwm|pwmList[9][9] .modeMux = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][9] .FeedbackMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][9] .ShiftMux = 1'b0;
defparam \macro_inst|controller|sm_pwm|pwmList[9][9] .BypassEn = 1'b1;
defparam \macro_inst|controller|sm_pwm|pwmList[9][9] .CarryEnb = 1'b0;

alta_slice \macro_inst|mem_ahb_hrdata[0]~0 (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [0]),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|mem_ahb_hrdata[0]~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|mem_ahb_hrdata[0]~0 .coord_x = 18;
defparam \macro_inst|mem_ahb_hrdata[0]~0 .coord_y = 11;
defparam \macro_inst|mem_ahb_hrdata[0]~0 .coord_z = 14;
defparam \macro_inst|mem_ahb_hrdata[0]~0 .mask = 16'hF000;
defparam \macro_inst|mem_ahb_hrdata[0]~0 .modeMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[0]~0 .FeedbackMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[0]~0 .ShiftMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[0]~0 .BypassEn = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[0]~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|mem_ahb_hrdata[12]~12 (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [12]),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|mem_ahb_hrdata[12]~12_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|mem_ahb_hrdata[12]~12 .coord_x = 14;
defparam \macro_inst|mem_ahb_hrdata[12]~12 .coord_y = 7;
defparam \macro_inst|mem_ahb_hrdata[12]~12 .coord_z = 14;
defparam \macro_inst|mem_ahb_hrdata[12]~12 .mask = 16'hF000;
defparam \macro_inst|mem_ahb_hrdata[12]~12 .modeMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[12]~12 .FeedbackMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[12]~12 .ShiftMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[12]~12 .BypassEn = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[12]~12 .CarryEnb = 1'b1;

alta_slice \macro_inst|mem_ahb_hrdata[13]~13 (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [13]),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|mem_ahb_hrdata[13]~13_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|mem_ahb_hrdata[13]~13 .coord_x = 17;
defparam \macro_inst|mem_ahb_hrdata[13]~13 .coord_y = 11;
defparam \macro_inst|mem_ahb_hrdata[13]~13 .coord_z = 15;
defparam \macro_inst|mem_ahb_hrdata[13]~13 .mask = 16'hF000;
defparam \macro_inst|mem_ahb_hrdata[13]~13 .modeMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[13]~13 .FeedbackMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[13]~13 .ShiftMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[13]~13 .BypassEn = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[13]~13 .CarryEnb = 1'b1;

alta_slice \macro_inst|mem_ahb_hrdata[17]~17 (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [17]),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|mem_ahb_hrdata[17]~17_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|mem_ahb_hrdata[17]~17 .coord_x = 14;
defparam \macro_inst|mem_ahb_hrdata[17]~17 .coord_y = 12;
defparam \macro_inst|mem_ahb_hrdata[17]~17 .coord_z = 2;
defparam \macro_inst|mem_ahb_hrdata[17]~17 .mask = 16'hF000;
defparam \macro_inst|mem_ahb_hrdata[17]~17 .modeMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[17]~17 .FeedbackMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[17]~17 .ShiftMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[17]~17 .BypassEn = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[17]~17 .CarryEnb = 1'b1;

alta_slice \macro_inst|mem_ahb_hrdata[18]~18 (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [18]),
	.C(vcc),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|mem_ahb_hrdata[18]~18_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|mem_ahb_hrdata[18]~18 .coord_x = 14;
defparam \macro_inst|mem_ahb_hrdata[18]~18 .coord_y = 11;
defparam \macro_inst|mem_ahb_hrdata[18]~18 .coord_z = 7;
defparam \macro_inst|mem_ahb_hrdata[18]~18 .mask = 16'hCC00;
defparam \macro_inst|mem_ahb_hrdata[18]~18 .modeMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[18]~18 .FeedbackMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[18]~18 .ShiftMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[18]~18 .BypassEn = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[18]~18 .CarryEnb = 1'b1;

alta_slice \macro_inst|mem_ahb_hrdata[21]~21 (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [21]),
	.C(vcc),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|mem_ahb_hrdata[21]~21_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|mem_ahb_hrdata[21]~21 .coord_x = 14;
defparam \macro_inst|mem_ahb_hrdata[21]~21 .coord_y = 7;
defparam \macro_inst|mem_ahb_hrdata[21]~21 .coord_z = 13;
defparam \macro_inst|mem_ahb_hrdata[21]~21 .mask = 16'hCC00;
defparam \macro_inst|mem_ahb_hrdata[21]~21 .modeMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[21]~21 .FeedbackMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[21]~21 .ShiftMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[21]~21 .BypassEn = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[21]~21 .CarryEnb = 1'b1;

alta_slice \macro_inst|mem_ahb_hrdata[25]~25 (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [25]),
	.C(vcc),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|mem_ahb_hrdata[25]~25_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|mem_ahb_hrdata[25]~25 .coord_x = 14;
defparam \macro_inst|mem_ahb_hrdata[25]~25 .coord_y = 7;
defparam \macro_inst|mem_ahb_hrdata[25]~25 .coord_z = 8;
defparam \macro_inst|mem_ahb_hrdata[25]~25 .mask = 16'hCC00;
defparam \macro_inst|mem_ahb_hrdata[25]~25 .modeMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[25]~25 .FeedbackMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[25]~25 .ShiftMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[25]~25 .BypassEn = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[25]~25 .CarryEnb = 1'b1;

alta_slice \macro_inst|mem_ahb_hrdata[5]~5 (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [5]),
	.C(vcc),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|mem_ahb_hrdata[5]~5_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|mem_ahb_hrdata[5]~5 .coord_x = 15;
defparam \macro_inst|mem_ahb_hrdata[5]~5 .coord_y = 11;
defparam \macro_inst|mem_ahb_hrdata[5]~5 .coord_z = 10;
defparam \macro_inst|mem_ahb_hrdata[5]~5 .mask = 16'hCC00;
defparam \macro_inst|mem_ahb_hrdata[5]~5 .modeMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[5]~5 .FeedbackMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[5]~5 .ShiftMux = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[5]~5 .BypassEn = 1'b0;
defparam \macro_inst|mem_ahb_hrdata[5]~5 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Add1~0 (
	.A(\macro_inst|serial_lim_input_inst|bit_counter [2]),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|bit_counter [1]),
	.D(\macro_inst|serial_lim_input_inst|bit_counter [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Add1~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Add1~0 .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|Add1~0 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|Add1~0 .coord_z = 10;
defparam \macro_inst|serial_lim_input_inst|Add1~0 .mask = 16'h5AAA;
defparam \macro_inst|serial_lim_input_inst|Add1~0 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Add1~0 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Add1~0 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Add1~0 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Add1~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Decoder0~0 (
	.A(\sys_resetn~clkctrl_outclk ),
	.B(\macro_inst|serial_lim_input_inst|shift_out_d~q ),
	.C(\macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT~q ),
	.D(\macro_inst|serial_lim_input_inst|shift_out~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Decoder0~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Decoder0~0 .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~0 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~0 .coord_z = 7;
defparam \macro_inst|serial_lim_input_inst|Decoder0~0 .mask = 16'h1000;
defparam \macro_inst|serial_lim_input_inst|Decoder0~0 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~0 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~0 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~0 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Decoder0~1 (
	.A(\macro_inst|serial_lim_input_inst|Decoder0~0_combout ),
	.B(\macro_inst|serial_lim_input_inst|bit_counter [0]),
	.C(\macro_inst|serial_lim_input_inst|bit_counter [1]),
	.D(\macro_inst|serial_lim_input_inst|bit_counter [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Decoder0~1_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Decoder0~1 .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|Decoder0~1 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~1 .coord_z = 1;
defparam \macro_inst|serial_lim_input_inst|Decoder0~1 .mask = 16'h2000;
defparam \macro_inst|serial_lim_input_inst|Decoder0~1 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~1 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~1 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~1 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~1 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Decoder0~2 (
	.A(\macro_inst|serial_lim_input_inst|bit_counter [2]),
	.B(\macro_inst|serial_lim_input_inst|bit_counter [1]),
	.C(\macro_inst|serial_lim_input_inst|bit_counter [0]),
	.D(\macro_inst|serial_lim_input_inst|Decoder0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Decoder0~2_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Decoder0~2 .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~2 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~2 .coord_z = 14;
defparam \macro_inst|serial_lim_input_inst|Decoder0~2 .mask = 16'h8000;
defparam \macro_inst|serial_lim_input_inst|Decoder0~2 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~2 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~2 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~2 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~2 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Decoder0~3 (
	.A(\macro_inst|serial_lim_input_inst|bit_counter [2]),
	.B(\macro_inst|serial_lim_input_inst|bit_counter [1]),
	.C(\macro_inst|serial_lim_input_inst|bit_counter [0]),
	.D(\macro_inst|serial_lim_input_inst|Decoder0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Decoder0~3_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Decoder0~3 .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~3 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~3 .coord_z = 10;
defparam \macro_inst|serial_lim_input_inst|Decoder0~3 .mask = 16'h0200;
defparam \macro_inst|serial_lim_input_inst|Decoder0~3 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~3 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~3 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~3 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~3 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Decoder0~4 (
	.A(\macro_inst|serial_lim_input_inst|bit_counter [1]),
	.B(\macro_inst|serial_lim_input_inst|bit_counter [0]),
	.C(\macro_inst|serial_lim_input_inst|bit_counter [2]),
	.D(\macro_inst|serial_lim_input_inst|Decoder0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Decoder0~4_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Decoder0~4 .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|Decoder0~4 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~4 .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|Decoder0~4 .mask = 16'h4000;
defparam \macro_inst|serial_lim_input_inst|Decoder0~4 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~4 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~4 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~4 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~4 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Decoder0~5 (
	.A(\macro_inst|serial_lim_input_inst|bit_counter [1]),
	.B(\macro_inst|serial_lim_input_inst|Decoder0~0_combout ),
	.C(\macro_inst|serial_lim_input_inst|bit_counter [2]),
	.D(\macro_inst|serial_lim_input_inst|bit_counter [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Decoder0~5_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Decoder0~5 .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|Decoder0~5 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~5 .coord_z = 7;
defparam \macro_inst|serial_lim_input_inst|Decoder0~5 .mask = 16'h0800;
defparam \macro_inst|serial_lim_input_inst|Decoder0~5 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~5 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~5 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~5 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~5 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Decoder0~6 (
	.A(\macro_inst|serial_lim_input_inst|bit_counter [0]),
	.B(\macro_inst|serial_lim_input_inst|bit_counter [1]),
	.C(\macro_inst|serial_lim_input_inst|bit_counter [2]),
	.D(\macro_inst|serial_lim_input_inst|Decoder0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Decoder0~6_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Decoder0~6 .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~6 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~6 .coord_z = 11;
defparam \macro_inst|serial_lim_input_inst|Decoder0~6 .mask = 16'h0400;
defparam \macro_inst|serial_lim_input_inst|Decoder0~6 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~6 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~6 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~6 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~6 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Decoder0~7 (
	.A(\macro_inst|serial_lim_input_inst|bit_counter [0]),
	.B(\macro_inst|serial_lim_input_inst|bit_counter [1]),
	.C(\macro_inst|serial_lim_input_inst|bit_counter [2]),
	.D(\macro_inst|serial_lim_input_inst|Decoder0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Decoder0~7_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Decoder0~7 .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~7 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~7 .coord_z = 12;
defparam \macro_inst|serial_lim_input_inst|Decoder0~7 .mask = 16'h0200;
defparam \macro_inst|serial_lim_input_inst|Decoder0~7 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~7 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~7 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~7 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~7 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Decoder0~8 (
	.A(\macro_inst|serial_lim_input_inst|bit_counter [0]),
	.B(\macro_inst|serial_lim_input_inst|bit_counter [1]),
	.C(\macro_inst|serial_lim_input_inst|bit_counter [2]),
	.D(\macro_inst|serial_lim_input_inst|Decoder0~0_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Decoder0~8_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Decoder0~8 .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~8 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|Decoder0~8 .coord_z = 1;
defparam \macro_inst|serial_lim_input_inst|Decoder0~8 .mask = 16'h0100;
defparam \macro_inst|serial_lim_input_inst|Decoder0~8 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~8 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~8 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~8 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Decoder0~8 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Equal0~0 (
	.A(\macro_inst|serial_lim_input_inst|load_counter [0]),
	.B(\macro_inst|serial_lim_input_inst|load_counter [1]),
	.C(\macro_inst|serial_lim_input_inst|load_counter [3]),
	.D(\macro_inst|serial_lim_input_inst|load_counter [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Equal0~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Equal0~0 .coord_x = 3;
defparam \macro_inst|serial_lim_input_inst|Equal0~0 .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|Equal0~0 .coord_z = 13;
defparam \macro_inst|serial_lim_input_inst|Equal0~0 .mask = 16'h0001;
defparam \macro_inst|serial_lim_input_inst|Equal0~0 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~0 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~0 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~0 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Equal0~1 (
	.A(\macro_inst|serial_lim_input_inst|load_counter [7]),
	.B(\macro_inst|serial_lim_input_inst|load_counter [4]),
	.C(\macro_inst|serial_lim_input_inst|load_counter [5]),
	.D(\macro_inst|serial_lim_input_inst|load_counter [6]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Equal0~1_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Equal0~1 .coord_x = 3;
defparam \macro_inst|serial_lim_input_inst|Equal0~1 .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|Equal0~1 .coord_z = 0;
defparam \macro_inst|serial_lim_input_inst|Equal0~1 .mask = 16'h0001;
defparam \macro_inst|serial_lim_input_inst|Equal0~1 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~1 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~1 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~1 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~1 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Equal0~2 (
	.A(\macro_inst|serial_lim_input_inst|load_counter [9]),
	.B(\macro_inst|serial_lim_input_inst|load_counter [10]),
	.C(\macro_inst|serial_lim_input_inst|load_counter [11]),
	.D(\macro_inst|serial_lim_input_inst|load_counter [8]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Equal0~2_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Equal0~2 .coord_x = 3;
defparam \macro_inst|serial_lim_input_inst|Equal0~2 .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|Equal0~2 .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|Equal0~2 .mask = 16'h0001;
defparam \macro_inst|serial_lim_input_inst|Equal0~2 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~2 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~2 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~2 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~2 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Equal0~3 (
	.A(\macro_inst|serial_lim_input_inst|load_counter [15]),
	.B(\macro_inst|serial_lim_input_inst|load_counter [13]),
	.C(\macro_inst|serial_lim_input_inst|load_counter [14]),
	.D(\macro_inst|serial_lim_input_inst|load_counter [12]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Equal0~3_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Equal0~3 .coord_x = 3;
defparam \macro_inst|serial_lim_input_inst|Equal0~3 .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|Equal0~3 .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|Equal0~3 .mask = 16'h0001;
defparam \macro_inst|serial_lim_input_inst|Equal0~3 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~3 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~3 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~3 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~3 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Equal0~4 (
	.A(\macro_inst|serial_lim_input_inst|Equal0~3_combout ),
	.B(\macro_inst|serial_lim_input_inst|Equal0~0_combout ),
	.C(\macro_inst|serial_lim_input_inst|Equal0~1_combout ),
	.D(\macro_inst|serial_lim_input_inst|Equal0~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Equal0~4_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Equal0~4 .coord_x = 3;
defparam \macro_inst|serial_lim_input_inst|Equal0~4 .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|Equal0~4 .coord_z = 4;
defparam \macro_inst|serial_lim_input_inst|Equal0~4 .mask = 16'h8000;
defparam \macro_inst|serial_lim_input_inst|Equal0~4 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~4 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~4 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~4 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal0~4 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Equal2~0 (
	.A(\macro_inst|serial_lim_input_inst|shift_div_counter [1]),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [3]),
	.C(\macro_inst|serial_lim_input_inst|shift_div_counter [0]),
	.D(\macro_inst|serial_lim_input_inst|shift_div_counter [2]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Equal2~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Equal2~0 .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|Equal2~0 .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|Equal2~0 .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|Equal2~0 .mask = 16'hFFBF;
defparam \macro_inst|serial_lim_input_inst|Equal2~0 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~0 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~0 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~0 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Equal2~1 (
	.A(\macro_inst|serial_lim_input_inst|shift_div_counter [6]),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [4]),
	.C(\macro_inst|serial_lim_input_inst|shift_div_counter [5]),
	.D(\macro_inst|serial_lim_input_inst|shift_div_counter [7]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Equal2~1_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Equal2~1 .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|Equal2~1 .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|Equal2~1 .coord_z = 6;
defparam \macro_inst|serial_lim_input_inst|Equal2~1 .mask = 16'hFFFE;
defparam \macro_inst|serial_lim_input_inst|Equal2~1 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~1 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~1 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~1 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~1 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Equal2~2 (
	.A(\macro_inst|serial_lim_input_inst|shift_div_counter [8]),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [11]),
	.C(\macro_inst|serial_lim_input_inst|shift_div_counter [10]),
	.D(\macro_inst|serial_lim_input_inst|shift_div_counter [9]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Equal2~2_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Equal2~2 .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|Equal2~2 .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|Equal2~2 .coord_z = 3;
defparam \macro_inst|serial_lim_input_inst|Equal2~2 .mask = 16'hFFFE;
defparam \macro_inst|serial_lim_input_inst|Equal2~2 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~2 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~2 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~2 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~2 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Equal2~3 (
	.A(\macro_inst|serial_lim_input_inst|shift_div_counter [14]),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [13]),
	.C(\macro_inst|serial_lim_input_inst|shift_div_counter [12]),
	.D(\macro_inst|serial_lim_input_inst|shift_div_counter [15]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Equal2~3_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Equal2~3 .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|Equal2~3 .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|Equal2~3 .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|Equal2~3 .mask = 16'hFFFE;
defparam \macro_inst|serial_lim_input_inst|Equal2~3 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~3 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~3 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~3 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~3 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Equal2~4 (
	.A(\macro_inst|serial_lim_input_inst|Equal2~3_combout ),
	.B(\macro_inst|serial_lim_input_inst|Equal2~0_combout ),
	.C(\macro_inst|serial_lim_input_inst|Equal2~1_combout ),
	.D(\macro_inst|serial_lim_input_inst|Equal2~2_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Equal2~4_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Equal2~4 .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|Equal2~4 .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|Equal2~4 .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|Equal2~4 .mask = 16'hFFFE;
defparam \macro_inst|serial_lim_input_inst|Equal2~4 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~4 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~4 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~4 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Equal2~4 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Selector20~2 (
	.A(\macro_inst|serial_lim_input_inst|Equal0~4_combout ),
	.B(\macro_inst|serial_lim_input_inst|shift_out_d~q ),
	.C(\macro_inst|serial_lim_input_inst|shift_out~q ),
	.D(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Selector20~2_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Selector20~2 .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|Selector20~2 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|Selector20~2 .coord_z = 11;
defparam \macro_inst|serial_lim_input_inst|Selector20~2 .mask = 16'h2000;
defparam \macro_inst|serial_lim_input_inst|Selector20~2 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Selector20~2 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Selector20~2 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Selector20~2 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Selector20~2 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Selector20~3 (
	.A(\macro_inst|serial_lim_input_inst|bit_counter [2]),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|bit_counter [1]),
	.D(\macro_inst|serial_lim_input_inst|bit_counter [0]),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Selector20~3_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Selector20~3 .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|Selector20~3 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|Selector20~3 .coord_z = 4;
defparam \macro_inst|serial_lim_input_inst|Selector20~3 .mask = 16'hA000;
defparam \macro_inst|serial_lim_input_inst|Selector20~3 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Selector20~3 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Selector20~3 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Selector20~3 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Selector20~3 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|Selector20~5 (
	.A(\macro_inst|serial_lim_input_inst|Selector20~3_combout ),
	.B(\macro_inst|serial_lim_input_inst|shift_out_d~q ),
	.C(\macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT~q ),
	.D(\macro_inst|serial_lim_input_inst|shift_out~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Selector20~5_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|Selector20~5 .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|Selector20~5 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|Selector20~5 .coord_z = 3;
defparam \macro_inst|serial_lim_input_inst|Selector20~5 .mask = 16'h2000;
defparam \macro_inst|serial_lim_input_inst|Selector20~5 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Selector20~5 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Selector20~5 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Selector20~5 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|Selector20~5 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|ahb_read_transfer (
	.A(\rv32.mem_ahb_hready ),
	.B(\rv32.mem_ahb_hwrite ),
	.C(\rv32.mem_ahb_htrans[1] ),
	.D(\macro_inst|Equal1~8_combout ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|ahb_read_transfer~combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|ahb_read_transfer .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|ahb_read_transfer .coord_y = 11;
defparam \macro_inst|serial_lim_input_inst|ahb_read_transfer .coord_z = 10;
defparam \macro_inst|serial_lim_input_inst|ahb_read_transfer .mask = 16'h2000;
defparam \macro_inst|serial_lim_input_inst|ahb_read_transfer .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|ahb_read_transfer .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|ahb_read_transfer .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|ahb_read_transfer .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|ahb_read_transfer .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|bit_counter[0] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|bit_counter[1]~1_combout ),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|bit_counter [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X46_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|bit_counter[0]~4_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|bit_counter [0]));
defparam \macro_inst|serial_lim_input_inst|bit_counter[0] .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|bit_counter[0] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|bit_counter[0] .coord_z = 6;
defparam \macro_inst|serial_lim_input_inst|bit_counter[0] .mask = 16'hC3C0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[0] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[0] .FeedbackMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|bit_counter[0] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[0] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[0] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|bit_counter[1] (
	.A(\macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT~q ),
	.B(\macro_inst|serial_lim_input_inst|bit_counter[1]~1_combout ),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|bit_counter [0]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|bit_counter [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X46_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|bit_counter[1]~3_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|bit_counter [1]));
defparam \macro_inst|serial_lim_input_inst|bit_counter[1] .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1] .coord_z = 8;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1] .mask = 16'hC2E0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1] .FeedbackMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|bit_counter[1]~0 (
	.A(\macro_inst|serial_lim_input_inst|Selector20~3_combout ),
	.B(\macro_inst|serial_lim_input_inst|shift_out_d~q ),
	.C(\macro_inst|serial_lim_input_inst|shift_out~q ),
	.D(\macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|bit_counter[1]~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~0 .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~0 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~0 .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~0 .mask = 16'hEFFF;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~0 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~0 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~0 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~0 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|bit_counter[1]~1 (
	.A(\macro_inst|serial_lim_input_inst|bit_counter[1]~0_combout ),
	.B(\macro_inst|serial_lim_input_inst|shift_rise~combout ),
	.C(\macro_inst|serial_lim_input_inst|Equal0~4_combout ),
	.D(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|bit_counter[1]~1_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~1 .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~1 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~1 .coord_z = 3;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~1 .mask = 16'h2AAA;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~1 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~1 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~1 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~1 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[1]~1 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|bit_counter[2] (
	.A(\macro_inst|serial_lim_input_inst|Add1~0_combout ),
	.B(\macro_inst|serial_lim_input_inst|bit_counter[1]~1_combout ),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|bit_counter [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X46_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|bit_counter[2]~2_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|bit_counter [2]));
defparam \macro_inst|serial_lim_input_inst|bit_counter[2] .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|bit_counter[2] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|bit_counter[2] .coord_z = 0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[2] .mask = 16'hE2C0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[2] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[2] .FeedbackMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|bit_counter[2] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[2] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|bit_counter[2] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|capture_done (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|Selector20~5_combout ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|capture_done~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X49_Y4_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|capture_done~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|capture_done~q ));
defparam \macro_inst|serial_lim_input_inst|capture_done .coord_x = 3;
defparam \macro_inst|serial_lim_input_inst|capture_done .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|capture_done .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|capture_done .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|capture_done .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|capture_done .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|capture_done .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|capture_done .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|capture_done .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[0][1]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X51_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[0]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [0]));
defparam \macro_inst|serial_lim_input_inst|captured_data[0] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[0] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[0] .coord_z = 11;
defparam \macro_inst|serial_lim_input_inst|captured_data[0] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[0] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[0] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[0] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[0] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[0] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[10] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|shift_buffer[1][3]~q ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [10]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[10]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [10]));
defparam \macro_inst|serial_lim_input_inst|captured_data[10] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[10] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[10] .coord_z = 1;
defparam \macro_inst|serial_lim_input_inst|captured_data[10] .mask = 16'hF0F0;
defparam \macro_inst|serial_lim_input_inst|captured_data[10] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[10] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[10] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[10] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[10] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[11] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[1][2]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [11]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[11]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [11]));
defparam \macro_inst|serial_lim_input_inst|captured_data[11] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[11] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[11] .coord_z = 12;
defparam \macro_inst|serial_lim_input_inst|captured_data[11] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[11] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[11] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[11] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[11] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[11] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[12] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[1][4]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [12]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[12]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [12]));
defparam \macro_inst|serial_lim_input_inst|captured_data[12] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[12] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[12] .coord_z = 3;
defparam \macro_inst|serial_lim_input_inst|captured_data[12] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[12] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[12] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[12] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[12] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[12] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[13] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|shift_buffer[1][5]~q ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [13]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[13]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [13]));
defparam \macro_inst|serial_lim_input_inst|captured_data[13] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[13] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[13] .coord_z = 3;
defparam \macro_inst|serial_lim_input_inst|captured_data[13] .mask = 16'hF0F0;
defparam \macro_inst|serial_lim_input_inst|captured_data[13] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[13] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[13] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[13] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[13] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[14] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[1][6]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [14]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[14]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [14]));
defparam \macro_inst|serial_lim_input_inst|captured_data[14] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[14] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[14] .coord_z = 14;
defparam \macro_inst|serial_lim_input_inst|captured_data[14] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[14] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[14] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[14] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[14] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[14] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[15] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[1][7]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [15]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[15]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [15]));
defparam \macro_inst|serial_lim_input_inst|captured_data[15] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[15] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[15] .coord_z = 11;
defparam \macro_inst|serial_lim_input_inst|captured_data[15] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[15] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[15] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[15] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[15] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[15] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[16] (
	.A(),
	.B(),
	.C(\macro_inst|serial_lim_input_inst|shift_buffer[2][1]~q ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [16]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X51_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y3_SIG ),
	.SyncReset(SyncReset_X51_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X51_Y3_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [16]));
defparam \macro_inst|serial_lim_input_inst|captured_data[16] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[16] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[16] .coord_z = 13;
defparam \macro_inst|serial_lim_input_inst|captured_data[16] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|captured_data[16] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|captured_data[16] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[16] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[16] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|captured_data[16] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[17] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[2][0]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [17]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X51_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[17]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [17]));
defparam \macro_inst|serial_lim_input_inst|captured_data[17] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[17] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[17] .coord_z = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[17] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[17] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[17] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[17] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[17] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[17] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[18] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_buffer[2][3]~q ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [18]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[18]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [18]));
defparam \macro_inst|serial_lim_input_inst|captured_data[18] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[18] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[18] .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|captured_data[18] .mask = 16'hCCCC;
defparam \macro_inst|serial_lim_input_inst|captured_data[18] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[18] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[18] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[18] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[18] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[19] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[2][2]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [19]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[19]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [19]));
defparam \macro_inst|serial_lim_input_inst|captured_data[19] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|captured_data[19] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[19] .coord_z = 3;
defparam \macro_inst|serial_lim_input_inst|captured_data[19] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[19] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[19] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[19] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[19] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[19] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[1] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[0][0]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[1]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [1]));
defparam \macro_inst|serial_lim_input_inst|captured_data[1] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[1] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[1] .coord_z = 6;
defparam \macro_inst|serial_lim_input_inst|captured_data[1] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[1] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[1] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[1] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[1] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[1] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[20] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[2][4]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [20]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X49_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[20]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [20]));
defparam \macro_inst|serial_lim_input_inst|captured_data[20] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[20] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|captured_data[20] .coord_z = 14;
defparam \macro_inst|serial_lim_input_inst|captured_data[20] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[20] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[20] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[20] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[20] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[20] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[21] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[2][5]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [21]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[21]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [21]));
defparam \macro_inst|serial_lim_input_inst|captured_data[21] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[21] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[21] .coord_z = 13;
defparam \macro_inst|serial_lim_input_inst|captured_data[21] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[21] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[21] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[21] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[21] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[21] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[22] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[2][6]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [22]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[22]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [22]));
defparam \macro_inst|serial_lim_input_inst|captured_data[22] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[22] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[22] .coord_z = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[22] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[22] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[22] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[22] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[22] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[22] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[23] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[2][7]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [23]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[23]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [23]));
defparam \macro_inst|serial_lim_input_inst|captured_data[23] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[23] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[23] .coord_z = 1;
defparam \macro_inst|serial_lim_input_inst|captured_data[23] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[23] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[23] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[23] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[23] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[23] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[24] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[3][1]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [24]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X51_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[24]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [24]));
defparam \macro_inst|serial_lim_input_inst|captured_data[24] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[24] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[24] .coord_z = 14;
defparam \macro_inst|serial_lim_input_inst|captured_data[24] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[24] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[24] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[24] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[24] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[24] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[25] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[3][0]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [25]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[25]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [25]));
defparam \macro_inst|serial_lim_input_inst|captured_data[25] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[25] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[25] .coord_z = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[25] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[25] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[25] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[25] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[25] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[25] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[26] (
	.A(\macro_inst|serial_lim_input_inst|shift_buffer[3][3]~q ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [26]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[26]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [26]));
defparam \macro_inst|serial_lim_input_inst|captured_data[26] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[26] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[26] .coord_z = 0;
defparam \macro_inst|serial_lim_input_inst|captured_data[26] .mask = 16'hAAAA;
defparam \macro_inst|serial_lim_input_inst|captured_data[26] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[26] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[26] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[26] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[26] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[27] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[3][2]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [27]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[27]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [27]));
defparam \macro_inst|serial_lim_input_inst|captured_data[27] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[27] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[27] .coord_z = 15;
defparam \macro_inst|serial_lim_input_inst|captured_data[27] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[27] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[27] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[27] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[27] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[27] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[28] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[3][4]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [28]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[28]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [28]));
defparam \macro_inst|serial_lim_input_inst|captured_data[28] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[28] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[28] .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|captured_data[28] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[28] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[28] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[28] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[28] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[28] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[29] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[3][5]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [29]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[29]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [29]));
defparam \macro_inst|serial_lim_input_inst|captured_data[29] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|captured_data[29] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[29] .coord_z = 1;
defparam \macro_inst|serial_lim_input_inst|captured_data[29] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[29] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[29] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[29] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[29] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[29] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[2] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[0][3]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[2]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [2]));
defparam \macro_inst|serial_lim_input_inst|captured_data[2] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[2] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[2] .coord_z = 6;
defparam \macro_inst|serial_lim_input_inst|captured_data[2] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[2] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[2] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[2] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[2] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[2] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[30] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[3][6]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [30]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[30]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [30]));
defparam \macro_inst|serial_lim_input_inst|captured_data[30] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|captured_data[30] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[30] .coord_z = 8;
defparam \macro_inst|serial_lim_input_inst|captured_data[30] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[30] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[30] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[30] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[30] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[30] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[31] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[3][7]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [31]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X51_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[31]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [31]));
defparam \macro_inst|serial_lim_input_inst|captured_data[31] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[31] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[31] .coord_z = 12;
defparam \macro_inst|serial_lim_input_inst|captured_data[31] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[31] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[31] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[31] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[31] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[31] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[32] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[4][1]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [32]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X51_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[32]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [32]));
defparam \macro_inst|serial_lim_input_inst|captured_data[32] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[32] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[32] .coord_z = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[32] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[32] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[32] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[32] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[32] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[32] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[33] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|shift_buffer[4][0]~q ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [33]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[33]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [33]));
defparam \macro_inst|serial_lim_input_inst|captured_data[33] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[33] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[33] .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|captured_data[33] .mask = 16'hF0F0;
defparam \macro_inst|serial_lim_input_inst|captured_data[33] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[33] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[33] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[33] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[33] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[34] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[4][3]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [34]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[34]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [34]));
defparam \macro_inst|serial_lim_input_inst|captured_data[34] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[34] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[34] .coord_z = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[34] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[34] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[34] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[34] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[34] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[34] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[35] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[4][2]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [35]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[35]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [35]));
defparam \macro_inst|serial_lim_input_inst|captured_data[35] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[35] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[35] .coord_z = 8;
defparam \macro_inst|serial_lim_input_inst|captured_data[35] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[35] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[35] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[35] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[35] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[35] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[36] (
	.A(),
	.B(),
	.C(\macro_inst|serial_lim_input_inst|shift_buffer[4][4]~q ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [36]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X49_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y2_SIG ),
	.SyncReset(SyncReset_X49_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X49_Y2_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [36]));
defparam \macro_inst|serial_lim_input_inst|captured_data[36] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[36] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|captured_data[36] .coord_z = 8;
defparam \macro_inst|serial_lim_input_inst|captured_data[36] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|captured_data[36] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|captured_data[36] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[36] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[36] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|captured_data[36] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[37] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[4][5]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [37]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[37]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [37]));
defparam \macro_inst|serial_lim_input_inst|captured_data[37] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|captured_data[37] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[37] .coord_z = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[37] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[37] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[37] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[37] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[37] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[37] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[38] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|shift_buffer[4][6]~q ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [38]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[38]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [38]));
defparam \macro_inst|serial_lim_input_inst|captured_data[38] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[38] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[38] .coord_z = 14;
defparam \macro_inst|serial_lim_input_inst|captured_data[38] .mask = 16'hF0F0;
defparam \macro_inst|serial_lim_input_inst|captured_data[38] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[38] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[38] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[38] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[38] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[39] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[4][7]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [39]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[39]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [39]));
defparam \macro_inst|serial_lim_input_inst|captured_data[39] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[39] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[39] .coord_z = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[39] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[39] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[39] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[39] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[39] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[39] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[3] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[0][2]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [3]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[3]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [3]));
defparam \macro_inst|serial_lim_input_inst|captured_data[3] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[3] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[3] .coord_z = 12;
defparam \macro_inst|serial_lim_input_inst|captured_data[3] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[3] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[3] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[3] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[3] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[3] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[40] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[5][1]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [40]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[40]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [40]));
defparam \macro_inst|serial_lim_input_inst|captured_data[40] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[40] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[40] .coord_z = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[40] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[40] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[40] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[40] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[40] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[40] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[41] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[5][0]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [41]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X51_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[41]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [41]));
defparam \macro_inst|serial_lim_input_inst|captured_data[41] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[41] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[41] .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|captured_data[41] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[41] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[41] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[41] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[41] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[41] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[42] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|shift_buffer[5][3]~q ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [42]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[42]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [42]));
defparam \macro_inst|serial_lim_input_inst|captured_data[42] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[42] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[42] .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[42] .mask = 16'hF0F0;
defparam \macro_inst|serial_lim_input_inst|captured_data[42] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[42] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[42] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[42] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[42] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[43] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[5][2]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [43]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[43]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [43]));
defparam \macro_inst|serial_lim_input_inst|captured_data[43] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[43] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[43] .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|captured_data[43] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[43] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[43] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[43] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[43] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[43] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[44] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[5][4]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [44]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X49_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y2_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[44]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [44]));
defparam \macro_inst|serial_lim_input_inst|captured_data[44] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[44] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|captured_data[44] .coord_z = 11;
defparam \macro_inst|serial_lim_input_inst|captured_data[44] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[44] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[44] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[44] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[44] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[44] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[45] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[5][5]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [45]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[45]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [45]));
defparam \macro_inst|serial_lim_input_inst|captured_data[45] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|captured_data[45] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[45] .coord_z = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[45] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[45] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[45] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[45] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[45] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[45] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[46] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[5][6]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [46]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[46]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [46]));
defparam \macro_inst|serial_lim_input_inst|captured_data[46] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|captured_data[46] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[46] .coord_z = 13;
defparam \macro_inst|serial_lim_input_inst|captured_data[46] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[46] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[46] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[46] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[46] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[46] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[47] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[5][7]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [47]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X53_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X53_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[47]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [47]));
defparam \macro_inst|serial_lim_input_inst|captured_data[47] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|captured_data[47] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[47] .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[47] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[47] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[47] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[47] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[47] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[47] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[4] (
	.A(),
	.B(),
	.C(\macro_inst|serial_lim_input_inst|shift_buffer[0][4]~q ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [4]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X49_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y2_SIG ),
	.SyncReset(SyncReset_X49_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X49_Y2_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [4]));
defparam \macro_inst|serial_lim_input_inst|captured_data[4] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[4] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|captured_data[4] .coord_z = 3;
defparam \macro_inst|serial_lim_input_inst|captured_data[4] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|captured_data[4] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|captured_data[4] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[4] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[4] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|captured_data[4] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[0][5]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [5]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[5]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [5]));
defparam \macro_inst|serial_lim_input_inst|captured_data[5] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|captured_data[5] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[5] .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|captured_data[5] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[5] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[5] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[5] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[5] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[5] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[6] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[0][6]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [6]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X49_Y4_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X49_Y4_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[6]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [6]));
defparam \macro_inst|serial_lim_input_inst|captured_data[6] .coord_x = 3;
defparam \macro_inst|serial_lim_input_inst|captured_data[6] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[6] .coord_z = 0;
defparam \macro_inst|serial_lim_input_inst|captured_data[6] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[6] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[6] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[6] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[6] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[6] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[7] (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|shift_buffer[0][7]~q ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [7]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[7]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [7]));
defparam \macro_inst|serial_lim_input_inst|captured_data[7] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[7] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[7] .coord_z = 13;
defparam \macro_inst|serial_lim_input_inst|captured_data[7] .mask = 16'hF0F0;
defparam \macro_inst|serial_lim_input_inst|captured_data[7] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[7] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[7] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[7] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[7] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[8] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_buffer[1][1]~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [8]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X51_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|captured_data[8]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [8]));
defparam \macro_inst|serial_lim_input_inst|captured_data[8] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[8] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[8] .coord_z = 10;
defparam \macro_inst|serial_lim_input_inst|captured_data[8] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|captured_data[8] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[8] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[8] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[8] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[8] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|captured_data[9] (
	.A(),
	.B(),
	.C(\macro_inst|serial_lim_input_inst|shift_buffer[1][0]~q ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|captured_data [9]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|capture_done~q_X51_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X51_Y3_SIG ),
	.SyncReset(SyncReset_X51_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X51_Y3_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|captured_data [9]));
defparam \macro_inst|serial_lim_input_inst|captured_data[9] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|captured_data[9] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|captured_data[9] .coord_z = 3;
defparam \macro_inst|serial_lim_input_inst|captured_data[9] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|captured_data[9] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|captured_data[9] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[9] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|captured_data[9] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|captured_data[9] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|load (
	.A(\macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT~q ),
	.B(\macro_inst|serial_lim_input_inst|load~0_combout ),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|Selector20~2_combout ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|load~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X47_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X47_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|load~1_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|load~q ));
defparam \macro_inst|serial_lim_input_inst|load .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|load .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|load .mask = 16'hA0E4;
defparam \macro_inst|serial_lim_input_inst|load .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load .FeedbackMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[0] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[0]~17_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[0]~18 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [0]));
defparam \macro_inst|serial_lim_input_inst|load_counter[0] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[0] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[0] .coord_z = 0;
defparam \macro_inst|serial_lim_input_inst|load_counter[0] .mask = 16'h33CC;
defparam \macro_inst|serial_lim_input_inst|load_counter[0] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[0] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[0] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[0] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[0] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[10] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [10]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[9]~37 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [10]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[10]~38_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[10]~39 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [10]));
defparam \macro_inst|serial_lim_input_inst|load_counter[10] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[10] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[10] .coord_z = 10;
defparam \macro_inst|serial_lim_input_inst|load_counter[10] .mask = 16'h3CCF;
defparam \macro_inst|serial_lim_input_inst|load_counter[10] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[10] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[10] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[10] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[10] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[11] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [11]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[10]~39 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [11]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[11]~40_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[11]~41 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [11]));
defparam \macro_inst|serial_lim_input_inst|load_counter[11] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[11] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[11] .coord_z = 11;
defparam \macro_inst|serial_lim_input_inst|load_counter[11] .mask = 16'hC303;
defparam \macro_inst|serial_lim_input_inst|load_counter[11] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[11] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[11] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[11] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[11] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[12] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [12]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[11]~41 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [12]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[12]~42_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[12]~43 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [12]));
defparam \macro_inst|serial_lim_input_inst|load_counter[12] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[12] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[12] .coord_z = 12;
defparam \macro_inst|serial_lim_input_inst|load_counter[12] .mask = 16'h3CCF;
defparam \macro_inst|serial_lim_input_inst|load_counter[12] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[12] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[12] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[12] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[12] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[13] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [13]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[12]~43 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [13]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[13]~44_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[13]~45 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [13]));
defparam \macro_inst|serial_lim_input_inst|load_counter[13] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[13] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[13] .coord_z = 13;
defparam \macro_inst|serial_lim_input_inst|load_counter[13] .mask = 16'hC303;
defparam \macro_inst|serial_lim_input_inst|load_counter[13] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[13] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[13] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[13] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[13] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[14] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [14]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[13]~45 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [14]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[14]~46_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[14]~47 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [14]));
defparam \macro_inst|serial_lim_input_inst|load_counter[14] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[14] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[14] .coord_z = 14;
defparam \macro_inst|serial_lim_input_inst|load_counter[14] .mask = 16'h3CCF;
defparam \macro_inst|serial_lim_input_inst|load_counter[14] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[14] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[14] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[14] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[14] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[14]~19 (
	.A(\macro_inst|serial_lim_input_inst|shift_rise~combout ),
	.B(\macro_inst|serial_lim_input_inst|load_counter[14]~16_combout ),
	.C(\macro_inst|serial_lim_input_inst|Equal0~4_combout ),
	.D(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[14]~19_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|load_counter[14]~19 .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[14]~19 .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|load_counter[14]~19 .coord_z = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[14]~19 .mask = 16'hCECC;
defparam \macro_inst|serial_lim_input_inst|load_counter[14]~19 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[14]~19 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[14]~19 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[14]~19 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[14]~19 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[15] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [15]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[14]~47 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [15]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[15]~48_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [15]));
defparam \macro_inst|serial_lim_input_inst|load_counter[15] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[15] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[15] .coord_z = 15;
defparam \macro_inst|serial_lim_input_inst|load_counter[15] .mask = 16'hC3C3;
defparam \macro_inst|serial_lim_input_inst|load_counter[15] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[15] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[15] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[15] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[15] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[1] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [1]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[0]~18 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[1]~20_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[1]~21 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [1]));
defparam \macro_inst|serial_lim_input_inst|load_counter[1] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[1] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[1] .coord_z = 1;
defparam \macro_inst|serial_lim_input_inst|load_counter[1] .mask = 16'hC303;
defparam \macro_inst|serial_lim_input_inst|load_counter[1] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[1] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[1] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[1] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[1] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[2] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [2]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[1]~21 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[2]~22_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[2]~23 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [2]));
defparam \macro_inst|serial_lim_input_inst|load_counter[2] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[2] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[2] .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|load_counter[2] .mask = 16'h3CCF;
defparam \macro_inst|serial_lim_input_inst|load_counter[2] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[2] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[2] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[2] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[2] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[3] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [3]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[2]~23 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [3]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[3]~24_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[3]~25 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [3]));
defparam \macro_inst|serial_lim_input_inst|load_counter[3] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[3] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[3] .coord_z = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[3] .mask = 16'hC303;
defparam \macro_inst|serial_lim_input_inst|load_counter[3] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[3] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[3] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[3] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[3] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[4] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [4]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[3]~25 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [4]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[4]~26_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[4]~27 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [4]));
defparam \macro_inst|serial_lim_input_inst|load_counter[4] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[4] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[4] .coord_z = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[4] .mask = 16'h3CCF;
defparam \macro_inst|serial_lim_input_inst|load_counter[4] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[4] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[4] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[4] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[4] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[5] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [5]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[4]~27 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [5]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[5]~28_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[5]~29 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [5]));
defparam \macro_inst|serial_lim_input_inst|load_counter[5] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[5] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[5] .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|load_counter[5] .mask = 16'hC303;
defparam \macro_inst|serial_lim_input_inst|load_counter[5] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[5] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[5] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[5] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[5] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[6] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [6]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[5]~29 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [6]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[6]~30_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[6]~31 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [6]));
defparam \macro_inst|serial_lim_input_inst|load_counter[6] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[6] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[6] .coord_z = 6;
defparam \macro_inst|serial_lim_input_inst|load_counter[6] .mask = 16'h3CCF;
defparam \macro_inst|serial_lim_input_inst|load_counter[6] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[6] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[6] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[6] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[6] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[7] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [7]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[6]~31 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [7]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[7]~32_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[7]~33 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [7]));
defparam \macro_inst|serial_lim_input_inst|load_counter[7] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[7] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[7] .coord_z = 7;
defparam \macro_inst|serial_lim_input_inst|load_counter[7] .mask = 16'hC303;
defparam \macro_inst|serial_lim_input_inst|load_counter[7] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[7] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[7] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[7] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[7] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[8] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [8]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[7]~33 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [8]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[8]~34_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[8]~35 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [8]));
defparam \macro_inst|serial_lim_input_inst|load_counter[8] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[8] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[8] .coord_z = 8;
defparam \macro_inst|serial_lim_input_inst|load_counter[8] .mask = 16'h3CCF;
defparam \macro_inst|serial_lim_input_inst|load_counter[8] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[8] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[8] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[8] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[8] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load_counter[9] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|load_counter [9]),
	.C(\~GND~combout ),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|load_counter[8]~35 ),
	.Qin(\macro_inst|serial_lim_input_inst|load_counter [9]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|load_counter[14]~19_combout_X46_Y2_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y2_SIG ),
	.SyncReset(SyncReset_X46_Y2_GND),
	.ShiftData(),
	.SyncLoad(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[9]~36_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|load_counter[9]~37 ),
	.Q(\macro_inst|serial_lim_input_inst|load_counter [9]));
defparam \macro_inst|serial_lim_input_inst|load_counter[9] .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load_counter[9] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|load_counter[9] .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|load_counter[9] .mask = 16'hC303;
defparam \macro_inst|serial_lim_input_inst|load_counter[9] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[9] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[9] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load_counter[9] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|load_counter[9] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|load~0 (
	.A(\macro_inst|serial_lim_input_inst|trigger_sync1~q ),
	.B(\macro_inst|serial_lim_input_inst|trigger_sync0~q ),
	.C(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q ),
	.D(\macro_inst|serial_lim_input_inst|load~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|load~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|load~0 .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|load~0 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|load~0 .coord_z = 13;
defparam \macro_inst|serial_lim_input_inst|load~0 .mask = 16'hF404;
defparam \macro_inst|serial_lim_input_inst|load~0 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load~0 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load~0 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load~0 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|load~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[0] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [32]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|serial_lim_input_inst|captured_data [0]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X56_Y5_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y5_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[0]~0_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [0]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[0] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[0] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[0] .coord_z = 11;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[0] .mask = 16'hCFC0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[0] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[0] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[0] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[0] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[0] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[10] (
	.A(\rv32.mem_ahb_haddr[2] ),
	.B(\macro_inst|serial_lim_input_inst|captured_data [10]),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|captured_data [42]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [10]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X56_Y5_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y5_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[10]~10_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [10]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[10] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[10] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[10] .coord_z = 0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[10] .mask = 16'hEE44;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[10] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[10] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[10] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[10] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[10] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[11] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [43]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|serial_lim_input_inst|captured_data [11]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [11]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X56_Y5_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y5_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[11]~11_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [11]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[11] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[11] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[11] .coord_z = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[11] .mask = 16'hCFC0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[11] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[11] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[11] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[11] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[11] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[12] (
	.A(\macro_inst|serial_lim_input_inst|captured_data [12]),
	.B(vcc),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|serial_lim_input_inst|captured_data [44]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [12]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X57_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y5_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X57_Y5_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y5_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[12]~12_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [12]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[12] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[12] .coord_y = 7;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[12] .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[12] .mask = 16'hFA0A;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[12] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[12] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[12] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[12] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[12] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[13] (
	.A(\macro_inst|serial_lim_input_inst|captured_data [45]),
	.B(vcc),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|serial_lim_input_inst|captured_data [13]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [13]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X56_Y3_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y3_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[13]~13_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [13]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[13] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[13] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[13] .coord_z = 0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[13] .mask = 16'hAFA0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[13] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[13] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[13] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[13] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[13] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[14] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [14]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|serial_lim_input_inst|captured_data [46]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [14]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X56_Y5_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y5_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[14]~14_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [14]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[14] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[14] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[14] .coord_z = 15;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[14] .mask = 16'hFC0C;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[14] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[14] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[14] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[14] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[14] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[15] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [47]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|serial_lim_input_inst|captured_data [15]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [15]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X57_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y5_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X57_Y5_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y5_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[15]~15_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [15]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[15] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[15] .coord_y = 7;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[15] .coord_z = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[15] .mask = 16'hCFC0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[15] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[15] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[15] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[15] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[15] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[16] (
	.A(\rv32.mem_ahb_haddr[2] ),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|captured_data [16]),
	.D(\rv32.mem_ahb_haddr[3] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [16]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[16]~16_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [16]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[16] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[16] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[16] .coord_z = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[16] .mask = 16'h0050;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[16] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[16] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[16] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[16] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[16] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[17] (
	.A(vcc),
	.B(\rv32.mem_ahb_haddr[3] ),
	.C(\macro_inst|serial_lim_input_inst|captured_data [17]),
	.D(\rv32.mem_ahb_haddr[2] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [17]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[17]~17_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [17]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[17] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[17] .coord_y = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[17] .coord_z = 8;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[17] .mask = 16'h0030;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[17] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[17] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[17] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[17] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[17] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[18] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [18]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\rv32.mem_ahb_haddr[3] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [18]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[18]~18_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [18]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[18] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[18] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[18] .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[18] .mask = 16'h000C;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[18] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[18] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[18] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[18] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[18] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[19] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [19]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\rv32.mem_ahb_haddr[3] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [19]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[19]~19_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [19]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[19] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[19] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[19] .coord_z = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[19] .mask = 16'h000C;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[19] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[19] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[19] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[19] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[19] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[1] (
	.A(\macro_inst|serial_lim_input_inst|captured_data [33]),
	.B(vcc),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|serial_lim_input_inst|captured_data [1]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X57_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y5_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X57_Y5_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y5_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[1]~1_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [1]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[1] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[1] .coord_y = 7;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[1] .coord_z = 3;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[1] .mask = 16'hAFA0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[1] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[1] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[1] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[1] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[1] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[20] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [20]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\rv32.mem_ahb_haddr[3] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [20]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[20]~20_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [20]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[20] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[20] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[20] .coord_z = 11;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[20] .mask = 16'h000C;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[20] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[20] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[20] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[20] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[20] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[21] (
	.A(\rv32.mem_ahb_haddr[2] ),
	.B(\rv32.mem_ahb_haddr[3] ),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|captured_data [21]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [21]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X57_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[21]~21_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [21]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[21] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[21] .coord_y = 7;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[21] .coord_z = 15;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[21] .mask = 16'h1100;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[21] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[21] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[21] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[21] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[21] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[22] (
	.A(vcc),
	.B(\rv32.mem_ahb_haddr[3] ),
	.C(\macro_inst|serial_lim_input_inst|captured_data [22]),
	.D(\rv32.mem_ahb_haddr[2] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [22]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[22]~22_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [22]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[22] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[22] .coord_y = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[22] .coord_z = 7;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[22] .mask = 16'h0030;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[22] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[22] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[22] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[22] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[22] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[23] (
	.A(\macro_inst|serial_lim_input_inst|captured_data [23]),
	.B(\rv32.mem_ahb_haddr[3] ),
	.C(vcc),
	.D(\rv32.mem_ahb_haddr[2] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [23]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[23]~23_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [23]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[23] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[23] .coord_y = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[23] .coord_z = 10;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[23] .mask = 16'h0022;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[23] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[23] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[23] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[23] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[23] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[24] (
	.A(vcc),
	.B(\rv32.mem_ahb_haddr[3] ),
	.C(\macro_inst|serial_lim_input_inst|captured_data [24]),
	.D(\rv32.mem_ahb_haddr[2] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [24]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[24]~24_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [24]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[24] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[24] .coord_y = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[24] .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[24] .mask = 16'h0030;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[24] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[24] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[24] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[24] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[24] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[25] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [25]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\rv32.mem_ahb_haddr[3] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [25]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X57_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y5_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[25]~25_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [25]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[25] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[25] .coord_y = 7;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[25] .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[25] .mask = 16'h000C;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[25] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[25] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[25] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[25] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[25] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[26] (
	.A(vcc),
	.B(\rv32.mem_ahb_haddr[3] ),
	.C(\macro_inst|serial_lim_input_inst|captured_data [26]),
	.D(\rv32.mem_ahb_haddr[2] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [26]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[26]~26_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [26]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[26] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[26] .coord_y = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[26] .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[26] .mask = 16'h0030;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[26] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[26] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[26] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[26] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[26] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[27] (
	.A(vcc),
	.B(\rv32.mem_ahb_haddr[2] ),
	.C(\macro_inst|serial_lim_input_inst|captured_data [27]),
	.D(\rv32.mem_ahb_haddr[3] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [27]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[27]~27_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [27]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[27] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[27] .coord_y = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[27] .coord_z = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[27] .mask = 16'h0030;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[27] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[27] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[27] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[27] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[27] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[28] (
	.A(vcc),
	.B(\rv32.mem_ahb_haddr[3] ),
	.C(\macro_inst|serial_lim_input_inst|captured_data [28]),
	.D(\rv32.mem_ahb_haddr[2] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [28]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X54_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X54_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[28]~28_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [28]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[28] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[28] .coord_y = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[28] .coord_z = 13;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[28] .mask = 16'h0030;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[28] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[28] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[28] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[28] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[28] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[29] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [29]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\rv32.mem_ahb_haddr[3] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [29]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[29]~29_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [29]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[29] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[29] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[29] .coord_z = 6;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[29] .mask = 16'h000C;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[29] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[29] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[29] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[29] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[29] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[2] (
	.A(\macro_inst|serial_lim_input_inst|captured_data [2]),
	.B(vcc),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|serial_lim_input_inst|captured_data [34]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X57_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y5_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X57_Y5_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y5_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[2]~2_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [2]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[2] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[2] .coord_y = 7;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[2] .coord_z = 10;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[2] .mask = 16'hFA0A;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[2] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[2] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[2] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[2] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[2] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[30] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [30]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\rv32.mem_ahb_haddr[3] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [30]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[30]~30_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [30]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[30] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[30] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[30] .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[30] .mask = 16'h000C;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[30] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[30] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[30] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[30] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[30] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[31] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [31]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\rv32.mem_ahb_haddr[3] ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [31]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[31]~31_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [31]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[31] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[31] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[31] .coord_z = 15;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[31] .mask = 16'h000C;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[31] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[31] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[31] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[31] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[31] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[3] (
	.A(\macro_inst|serial_lim_input_inst|captured_data [35]),
	.B(\macro_inst|serial_lim_input_inst|captured_data [3]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [3]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X57_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y5_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X57_Y5_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y5_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[3]~3_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [3]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[3] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[3] .coord_y = 7;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[3] .coord_z = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[3] .mask = 16'hACAC;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[3] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[3] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[3] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[3] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[3] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[4] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [36]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|serial_lim_input_inst|captured_data [4]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [4]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X57_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y5_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X57_Y5_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y5_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[4]~4_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [4]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[4] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[4] .coord_y = 7;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[4] .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[4] .mask = 16'hCFC0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[4] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[4] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[4] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[4] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[4] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[5] (
	.A(\macro_inst|serial_lim_input_inst|captured_data [5]),
	.B(vcc),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|serial_lim_input_inst|captured_data [37]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [5]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y3_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y3_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X56_Y3_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y3_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[5]~5_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [5]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[5] .coord_x = 12;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[5] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[5] .coord_z = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[5] .mask = 16'hFA0A;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[5] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[5] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[5] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[5] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[5] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[6] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [38]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|serial_lim_input_inst|captured_data [6]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [6]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X57_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y5_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X57_Y5_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y5_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[6]~6_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [6]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[6] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[6] .coord_y = 7;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[6] .coord_z = 6;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[6] .mask = 16'hCFC0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[6] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[6] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[6] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[6] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[6] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[7] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [39]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|serial_lim_input_inst|captured_data [7]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [7]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X57_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y5_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X57_Y5_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y5_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[7]~7_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [7]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[7] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[7] .coord_y = 7;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[7] .coord_z = 7;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[7] .mask = 16'hCFC0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[7] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[7] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[7] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[7] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[7] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[8] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|captured_data [8]),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|serial_lim_input_inst|captured_data [40]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [8]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X57_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X57_Y5_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X57_Y5_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X57_Y5_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[8]~8_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [8]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[8] .coord_x = 14;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[8] .coord_y = 7;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[8] .coord_z = 11;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[8] .mask = 16'hFC0C;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[8] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[8] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[8] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[8] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[8] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[9] (
	.A(\macro_inst|serial_lim_input_inst|captured_data [41]),
	.B(vcc),
	.C(\rv32.mem_ahb_haddr[2] ),
	.D(\macro_inst|serial_lim_input_inst|captured_data [9]),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [9]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|ahb_read_transfer~combout_X56_Y5_SIG_SIG ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X56_Y5_SIG ),
	.SyncReset(\rv32.mem_ahb_haddr[3]__SyncReset_X56_Y5_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X56_Y5_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|read_chunk[9]~9_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|mem_ahb_hrdata [9]));
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[9] .coord_x = 10;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[9] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[9] .coord_z = 8;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[9] .mask = 16'hAFA0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[9] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[9] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[9] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[9] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|mem_ahb_hrdata[9] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift (
	.A(vcc),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|load~q ),
	.D(\macro_inst|serial_lim_input_inst|shift_out~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift~combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|shift .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|shift .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift .coord_z = 4;
defparam \macro_inst|serial_lim_input_inst|shift .mask = 16'h0F00;
defparam \macro_inst|serial_lim_input_inst|shift .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[0][0] (
	.A(vcc),
	.B(vcc),
	.C(\LM_D0~input_o ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[0][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~2_combout_X51_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X51_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[0][0]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[0][0]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][0] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][0] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][0] .coord_z = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][0] .mask = 16'hF0F0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][0] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][0] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][0] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][0] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[0][1] (
	.A(\LM_D0~input_o ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[0][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~1_combout_X50_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X50_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[0][1]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[0][1]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][1] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][1] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][1] .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][1] .mask = 16'hAAAA;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][1] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][1] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][1] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][1] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][1] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[0][2] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D0~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[0][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~4_combout_X49_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[0][2]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[0][2]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][2] .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][2] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][2] .coord_z = 13;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][2] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][2] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][2] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][2] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][2] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][2] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[0][3] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D0~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[0][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~3_combout_X52_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X52_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[0][3]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[0][3]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][3] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][3] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][3] .coord_z = 11;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][3] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][3] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][3] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][3] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][3] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][3] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[0][4] (
	.A(),
	.B(),
	.C(\LM_D0~input_o ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[0][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~5_combout_X49_Y2_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y2_GND),
	.SyncReset(SyncReset_X49_Y2_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X49_Y2_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[0][4]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][4] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][4] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][4] .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][4] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][4] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][4] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][4] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][4] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][4] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[0][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D0~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[0][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~6_combout_X52_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X52_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[0][5]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[0][5]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][5] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][5] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][5] .coord_z = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][5] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][5] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][5] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][5] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][5] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[0][6] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D0~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[0][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~7_combout_X49_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[0][6]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[0][6]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][6] .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][6] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][6] .coord_z = 12;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][6] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][6] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][6] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][6] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][6] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[0][7] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D0~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[0][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~8_combout_X50_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X50_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[0][7]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[0][7]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][7] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][7] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][7] .coord_z = 12;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][7] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][7] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][7] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][7] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][7] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[0][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[1][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D1~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[1][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~2_combout_X51_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X51_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[1][0]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[1][0]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][0] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][0] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][0] .coord_z = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][0] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][0] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][0] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][0] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][0] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[1][1] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D1~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[1][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~1_combout_X50_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X50_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[1][1]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[1][1]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][1] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][1] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][1] .coord_z = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][1] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][1] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][1] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][1] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][1] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][1] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[1][2] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D1~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[1][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~4_combout_X49_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[1][2]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[1][2]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][2] .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][2] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][2] .coord_z = 11;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][2] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][2] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][2] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][2] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][2] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][2] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[1][3] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D1~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[1][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~3_combout_X52_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X52_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[1][3]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[1][3]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][3] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][3] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][3] .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][3] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][3] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][3] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][3] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][3] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][3] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[1][4] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D1~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[1][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~5_combout_X49_Y2_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y2_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[1][4]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[1][4]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][4] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][4] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][4] .coord_z = 12;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][4] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][4] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][4] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][4] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][4] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][4] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[1][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D1~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[1][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~6_combout_X52_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X52_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[1][5]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[1][5]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][5] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][5] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][5] .coord_z = 15;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][5] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][5] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][5] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][5] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][5] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[1][6] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D1~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[1][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~7_combout_X49_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[1][6]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[1][6]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][6] .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][6] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][6] .coord_z = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][6] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][6] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][6] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][6] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][6] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[1][7] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D1~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[1][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~8_combout_X50_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X50_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[1][7]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[1][7]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][7] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][7] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][7] .coord_z = 11;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][7] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][7] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][7] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][7] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][7] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[1][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[2][0] (
	.A(),
	.B(),
	.C(\LM_D2~input_o ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[2][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~2_combout_X51_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X51_Y3_GND),
	.SyncReset(SyncReset_X51_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X51_Y3_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[2][0]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][0] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][0] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][0] .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][0] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][0] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][0] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][0] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][0] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[2][1] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D2~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[2][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~1_combout_X50_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X50_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[2][1]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[2][1]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][1] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][1] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][1] .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][1] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][1] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][1] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][1] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][1] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][1] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[2][2] (
	.A(),
	.B(),
	.C(\LM_D2~input_o ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[2][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~4_combout_X49_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y3_GND),
	.SyncReset(SyncReset_X49_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X49_Y3_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[2][2]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][2] .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][2] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][2] .coord_z = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][2] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][2] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][2] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][2] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][2] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][2] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[2][3] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D2~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[2][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~3_combout_X52_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X52_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[2][3]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[2][3]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][3] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][3] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][3] .coord_z = 10;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][3] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][3] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][3] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][3] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][3] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][3] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[2][4] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D2~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[2][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~5_combout_X49_Y2_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y2_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[2][4]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[2][4]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][4] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][4] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][4] .coord_z = 1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][4] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][4] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][4] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][4] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][4] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][4] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[2][5] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D2~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[2][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~6_combout_X52_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X52_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[2][5]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[2][5]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][5] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][5] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][5] .coord_z = 7;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][5] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][5] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][5] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][5] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][5] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[2][6] (
	.A(),
	.B(),
	.C(\LM_D2~input_o ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[2][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~7_combout_X49_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y3_GND),
	.SyncReset(SyncReset_X49_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X49_Y3_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[2][6]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][6] .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][6] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][6] .coord_z = 1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][6] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][6] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][6] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][6] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][6] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[2][7] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D2~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[2][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~8_combout_X50_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X50_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[2][7]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[2][7]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][7] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][7] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][7] .coord_z = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][7] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][7] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][7] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][7] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][7] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[2][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[3][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D3~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[3][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~2_combout_X51_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X51_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[3][0]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[3][0]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][0] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][0] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][0] .coord_z = 0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][0] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][0] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][0] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][0] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][0] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[3][1] (
	.A(),
	.B(),
	.C(\LM_D3~input_o ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[3][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~1_combout_X50_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X50_Y3_GND),
	.SyncReset(SyncReset_X50_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X50_Y3_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[3][1]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][1] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][1] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][1] .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][1] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][1] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][1] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][1] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][1] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][1] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[3][2] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D3~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[3][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~4_combout_X49_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[3][2]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[3][2]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][2] .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][2] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][2] .coord_z = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][2] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][2] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][2] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][2] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][2] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][2] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[3][3] (
	.A(),
	.B(),
	.C(\LM_D3~input_o ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[3][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~3_combout_X52_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X52_Y3_GND),
	.SyncReset(SyncReset_X52_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X52_Y3_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[3][3]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][3] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][3] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][3] .coord_z = 13;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][3] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][3] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][3] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][3] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][3] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][3] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[3][4] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D3~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[3][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~5_combout_X49_Y2_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y2_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[3][4]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[3][4]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][4] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][4] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][4] .coord_z = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][4] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][4] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][4] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][4] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][4] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][4] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[3][5] (
	.A(),
	.B(),
	.C(\LM_D3~input_o ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[3][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~6_combout_X52_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X52_Y3_GND),
	.SyncReset(SyncReset_X52_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X52_Y3_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[3][5]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][5] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][5] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][5] .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][5] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][5] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][5] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][5] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][5] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[3][6] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D3~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[3][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~7_combout_X49_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[3][6]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[3][6]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][6] .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][6] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][6] .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][6] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][6] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][6] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][6] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][6] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[3][7] (
	.A(),
	.B(),
	.C(\LM_D3~input_o ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[3][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~8_combout_X50_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X50_Y3_GND),
	.SyncReset(SyncReset_X50_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X50_Y3_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[3][7]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][7] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][7] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][7] .coord_z = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][7] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][7] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][7] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][7] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][7] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[3][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[4][0] (
	.A(),
	.B(),
	.C(\LM_D4~input_o ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[4][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~2_combout_X51_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X51_Y3_GND),
	.SyncReset(SyncReset_X51_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X51_Y3_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[4][0]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][0] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][0] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][0] .coord_z = 15;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][0] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][0] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][0] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][0] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][0] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[4][1] (
	.A(vcc),
	.B(vcc),
	.C(\LM_D4~input_o ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[4][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~1_combout_X50_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X50_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[4][1]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[4][1]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][1] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][1] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][1] .coord_z = 7;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][1] .mask = 16'hF0F0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][1] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][1] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][1] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][1] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][1] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[4][2] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D4~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[4][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~4_combout_X49_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[4][2]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[4][2]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][2] .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][2] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][2] .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][2] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][2] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][2] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][2] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][2] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][2] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[4][3] (
	.A(\LM_D4~input_o ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[4][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~3_combout_X52_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X52_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[4][3]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[4][3]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][3] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][3] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][3] .coord_z = 14;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][3] .mask = 16'hAAAA;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][3] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][3] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][3] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][3] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][3] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[4][4] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D4~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[4][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~5_combout_X49_Y2_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y2_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[4][4]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[4][4]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][4] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][4] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][4] .coord_z = 0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][4] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][4] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][4] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][4] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][4] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][4] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[4][5] (
	.A(\LM_D4~input_o ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[4][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~6_combout_X52_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X52_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[4][5]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[4][5]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][5] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][5] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][5] .coord_z = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][5] .mask = 16'hAAAA;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][5] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][5] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][5] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][5] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[4][6] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D4~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[4][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~7_combout_X49_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[4][6]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[4][6]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][6] .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][6] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][6] .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][6] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][6] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][6] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][6] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][6] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[4][7] (
	.A(vcc),
	.B(vcc),
	.C(\LM_D4~input_o ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[4][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~8_combout_X50_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X50_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[4][7]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[4][7]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][7] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][7] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][7] .coord_z = 14;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][7] .mask = 16'hF0F0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][7] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][7] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][7] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][7] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[4][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[5][0] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D5~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[5][0]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~2_combout_X51_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X51_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[5][0]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[5][0]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][0] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][0] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][0] .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][0] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][0] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][0] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][0] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][0] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][0] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[5][1] (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\LM_D5~input_o ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[5][1]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~1_combout_X50_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X50_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[5][1]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[5][1]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][1] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][1] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][1] .coord_z = 13;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][1] .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][1] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][1] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][1] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][1] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][1] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[5][2] (
	.A(),
	.B(),
	.C(\LM_D5~input_o ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[5][2]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~4_combout_X49_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y3_GND),
	.SyncReset(SyncReset_X49_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X49_Y3_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[5][2]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][2] .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][2] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][2] .coord_z = 10;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][2] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][2] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][2] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][2] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][2] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][2] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[5][3] (
	.A(\LM_D5~input_o ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[5][3]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~3_combout_X52_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X52_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[5][3]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[5][3]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][3] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][3] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][3] .coord_z = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][3] .mask = 16'hAAAA;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][3] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][3] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][3] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][3] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][3] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[5][4] (
	.A(vcc),
	.B(vcc),
	.C(\LM_D5~input_o ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[5][4]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~5_combout_X49_Y2_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y2_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[5][4]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[5][4]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][4] .coord_x = 9;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][4] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][4] .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][4] .mask = 16'hF0F0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][4] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][4] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][4] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][4] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][4] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[5][5] (
	.A(\LM_D5~input_o ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[5][5]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~6_combout_X52_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X52_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[5][5]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[5][5]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][5] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][5] .coord_y = 3;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][5] .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][5] .mask = 16'hAAAA;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][5] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][5] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][5] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][5] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][5] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[5][6] (
	.A(),
	.B(),
	.C(\LM_D5~input_o ),
	.D(),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[5][6]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~7_combout_X49_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X49_Y3_GND),
	.SyncReset(SyncReset_X49_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X49_Y3_VCC),
	.LutOut(),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[5][6]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][6] .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][6] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][6] .coord_z = 0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][6] .mask = 16'hFFFF;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][6] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][6] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][6] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][6] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][6] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_buffer[5][7] (
	.A(\LM_D5~input_o ),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_buffer[5][7]~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp__macro_inst|serial_lim_input_inst|Decoder0~8_combout_X50_Y3_SIG_SIG ),
	.AsyncReset(AsyncReset_X50_Y3_GND),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_buffer[5][7]~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_buffer[5][7]~q ));
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][7] .coord_x = 8;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][7] .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][7] .coord_z = 10;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][7] .mask = 16'hAAAA;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][7] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][7] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][7] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][7] .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_buffer[5][7] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[0] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [0]),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [0]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[0]~16_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[0]~17 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [0]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[0] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[0] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[0] .coord_z = 0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[0] .mask = 16'h33CC;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[0] .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[0] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[0] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[0] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[0] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[10] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [10]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[9]~36 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [10]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[10]~37_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[10]~38 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [10]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[10] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[10] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[10] .coord_z = 10;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[10] .mask = 16'hC30C;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[10] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[10] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[10] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[10] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[10] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[11] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [11]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[10]~38 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [11]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[11]~39_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[11]~40 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [11]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[11] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[11] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[11] .coord_z = 11;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[11] .mask = 16'h3C3F;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[11] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[11] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[11] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[11] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[11] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[12] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [12]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[11]~40 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [12]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[12]~41_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[12]~42 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [12]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[12] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[12] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[12] .coord_z = 12;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[12] .mask = 16'hC30C;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[12] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[12] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[12] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[12] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[12] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[13] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [13]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[12]~42 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [13]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[13]~43_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[13]~44 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [13]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[13] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[13] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[13] .coord_z = 13;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[13] .mask = 16'h3C3F;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[13] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[13] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[13] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[13] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[13] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[14] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [14]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[13]~44 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [14]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[14]~45_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[14]~46 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [14]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[14] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[14] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[14] .coord_z = 14;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[14] .mask = 16'hC30C;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[14] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[14] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[14] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[14] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[14] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[15] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [15]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[14]~46 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [15]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[15]~47_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [15]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[15] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[15] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[15] .coord_z = 15;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[15] .mask = 16'h3C3C;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[15] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[15] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[15] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[15] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[15] .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[1] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [1]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[0]~17 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [1]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[1]~18_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[1]~19 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [1]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[1] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[1] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[1] .coord_z = 1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[1] .mask = 16'h3C3F;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[1] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[1] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[1] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[1] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[1] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[2] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [2]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[1]~19 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [2]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~21_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~22 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [2]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2] .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2] .mask = 16'hC30C;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[2]~20 (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|Equal2~4_combout ),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|shift_enable~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2]~20 .coord_x = 6;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2]~20 .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2]~20 .coord_z = 0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2]~20 .mask = 16'h33FF;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2]~20 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2]~20 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2]~20 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2]~20 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[2]~20 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[3] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [3]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~22 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [3]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[3]~23_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[3]~24 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [3]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[3] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[3] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[3] .coord_z = 3;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[3] .mask = 16'h3C3F;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[3] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[3] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[3] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[3] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[3] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[4] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [4]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[3]~24 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [4]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[4]~25_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[4]~26 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [4]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[4] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[4] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[4] .coord_z = 4;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[4] .mask = 16'hC30C;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[4] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[4] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[4] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[4] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[4] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[5] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [5]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[4]~26 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [5]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[5]~27_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[5]~28 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [5]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[5] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[5] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[5] .coord_z = 5;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[5] .mask = 16'h3C3F;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[5] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[5] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[5] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[5] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[5] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[6] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [6]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[5]~28 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [6]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[6]~29_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[6]~30 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [6]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[6] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[6] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[6] .coord_z = 6;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[6] .mask = 16'hC30C;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[6] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[6] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[6] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[6] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[6] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[7] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [7]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[6]~30 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [7]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[7]~31_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[7]~32 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [7]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[7] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[7] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[7] .coord_z = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[7] .mask = 16'h3C3F;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[7] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[7] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[7] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[7] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[7] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[8] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [8]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[7]~32 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [8]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[8]~33_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[8]~34 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [8]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[8] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[8] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[8] .coord_z = 8;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[8] .mask = 16'hC30C;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[8] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[8] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[8] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[8] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[8] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_div_counter[9] (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_div_counter [9]),
	.C(vcc),
	.D(vcc),
	.Cin(\macro_inst|serial_lim_input_inst|shift_div_counter[8]~34 ),
	.Qin(\macro_inst|serial_lim_input_inst|shift_div_counter [9]),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X43_Y2_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X43_Y2_SIG ),
	.SyncReset(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ),
	.ShiftData(),
	.SyncLoad(SyncLoad_X43_Y2_GND),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_div_counter[9]~35_combout ),
	.Cout(\macro_inst|serial_lim_input_inst|shift_div_counter[9]~36 ),
	.Q(\macro_inst|serial_lim_input_inst|shift_div_counter [9]));
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[9] .coord_x = 7;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[9] .coord_y = 2;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[9] .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[9] .mask = 16'h3C3F;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[9] .modeMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[9] .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[9] .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[9] .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_div_counter[9] .CarryEnb = 1'b0;

alta_slice \macro_inst|serial_lim_input_inst|shift_enable (
	.A(vcc),
	.B(\macro_inst|serial_lim_input_inst|shift_enable~1_combout ),
	.C(\macro_inst|serial_lim_input_inst|shift_enable~0_combout ),
	.D(\macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_enable~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X46_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_enable~2_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_enable~q ));
defparam \macro_inst|serial_lim_input_inst|shift_enable .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|shift_enable .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_enable .coord_z = 12;
defparam \macro_inst|serial_lim_input_inst|shift_enable .mask = 16'hF0FC;
defparam \macro_inst|serial_lim_input_inst|shift_enable .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_enable .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_enable .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_enable .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_enable .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_enable~0 (
	.A(\macro_inst|serial_lim_input_inst|Selector20~3_combout ),
	.B(\macro_inst|serial_lim_input_inst|shift_rise~combout ),
	.C(\macro_inst|serial_lim_input_inst|shift_enable~q ),
	.D(\macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_enable~0_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|shift_enable~0 .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|shift_enable~0 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_enable~0 .coord_z = 13;
defparam \macro_inst|serial_lim_input_inst|shift_enable~0 .mask = 16'h7000;
defparam \macro_inst|serial_lim_input_inst|shift_enable~0 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_enable~0 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_enable~0 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_enable~0 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_enable~0 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_enable~1 (
	.A(\macro_inst|serial_lim_input_inst|shift_enable~q ),
	.B(\macro_inst|serial_lim_input_inst|trigger_sync0~q ),
	.C(\macro_inst|serial_lim_input_inst|trigger_sync1~q ),
	.D(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q ),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_enable~1_combout ),
	.Cout(),
	.Q());
defparam \macro_inst|serial_lim_input_inst|shift_enable~1 .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|shift_enable~1 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_enable~1 .coord_z = 15;
defparam \macro_inst|serial_lim_input_inst|shift_enable~1 .mask = 16'hAA0C;
defparam \macro_inst|serial_lim_input_inst|shift_enable~1 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_enable~1 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_enable~1 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_enable~1 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_enable~1 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_out (
	.A(\macro_inst|serial_lim_input_inst|shift_enable~q ),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|Equal2~4_combout ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_out~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X46_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_out~0_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_out~q ));
defparam \macro_inst|serial_lim_input_inst|shift_out .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|shift_out .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_out .coord_z = 14;
defparam \macro_inst|serial_lim_input_inst|shift_out .mask = 16'hA00A;
defparam \macro_inst|serial_lim_input_inst|shift_out .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_out .FeedbackMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_out .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_out .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_out .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|shift_out_d (
	.A(\macro_inst|serial_lim_input_inst|shift_out~q ),
	.B(vcc),
	.C(\macro_inst|serial_lim_input_inst|shift_out~q ),
	.D(vcc),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|shift_out_d~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X46_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X46_Y3_SIG ),
	.SyncReset(SyncReset_X46_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X46_Y3_VCC),
	.LutOut(\macro_inst|serial_lim_input_inst|shift_rise~combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|shift_out_d~q ));
defparam \macro_inst|serial_lim_input_inst|shift_out_d .coord_x = 5;
defparam \macro_inst|serial_lim_input_inst|shift_out_d .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|shift_out_d .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|shift_out_d .mask = 16'h0A0A;
defparam \macro_inst|serial_lim_input_inst|shift_out_d .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_out_d .FeedbackMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_out_d .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|shift_out_d .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|shift_out_d .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|state_reg.STATE_IDLE (
	.A(\macro_inst|serial_lim_input_inst|trigger_sync1~q ),
	.B(\macro_inst|serial_lim_input_inst|Selector20~5_combout ),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|trigger_sync0~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|state_reg.STATE_IDLE~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X47_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X47_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Selector18~0_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|state_reg.STATE_IDLE~q ));
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_IDLE .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_IDLE .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_IDLE .coord_z = 8;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_IDLE .mask = 16'h3130;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_IDLE .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_IDLE .FeedbackMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_IDLE .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_IDLE .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_IDLE .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD (
	.A(\macro_inst|serial_lim_input_inst|Selector20~5_combout ),
	.B(\macro_inst|serial_lim_input_inst|load_counter[14]~16_combout ),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|Selector20~2_combout ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X47_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X47_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Selector19~0_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q ));
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD .coord_z = 2;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD .mask = 16'h0054;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD .FeedbackMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT (
	.A(\macro_inst|serial_lim_input_inst|Selector20~5_combout ),
	.B(\macro_inst|serial_lim_input_inst|Selector20~2_combout ),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|load_counter[14]~16_combout ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X47_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X47_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|Selector20~4_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT~q ));
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT .coord_z = 6;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT .mask = 16'h4454;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT .FeedbackMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|state_reg.STATE_SHIFT .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|trigger_sync0 (
	.A(\macro_inst|serial_lim_input_inst|trigger_sync1~q ),
	.B(vcc),
	.C(\macro_inst|clock10Hz~q ),
	.D(\macro_inst|serial_lim_input_inst|state_reg.STATE_IDLE~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|trigger_sync0~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X47_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X47_Y3_SIG ),
	.SyncReset(SyncReset_X47_Y3_GND),
	.ShiftData(),
	.SyncLoad(SyncLoad_X47_Y3_VCC),
	.LutOut(\macro_inst|serial_lim_input_inst|load_counter[14]~16_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|trigger_sync0~q ));
defparam \macro_inst|serial_lim_input_inst|trigger_sync0 .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|trigger_sync0 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|trigger_sync0 .coord_z = 9;
defparam \macro_inst|serial_lim_input_inst|trigger_sync0 .mask = 16'h0050;
defparam \macro_inst|serial_lim_input_inst|trigger_sync0 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|trigger_sync0 .FeedbackMux = 1'b1;
defparam \macro_inst|serial_lim_input_inst|trigger_sync0 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|trigger_sync0 .BypassEn = 1'b1;
defparam \macro_inst|serial_lim_input_inst|trigger_sync0 .CarryEnb = 1'b1;

alta_slice \macro_inst|serial_lim_input_inst|trigger_sync1 (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(\macro_inst|serial_lim_input_inst|trigger_sync0~q ),
	.Cin(),
	.Qin(\macro_inst|serial_lim_input_inst|trigger_sync1~q ),
	.Clk(\auto_generated_inst.hbo_22_f9ff3d300b43c0f2_bp_X47_Y3_SIG_VCC ),
	.AsyncReset(\sys_resetn~clkctrl_outclk__AsyncReset_X47_Y3_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\macro_inst|serial_lim_input_inst|trigger_sync1~feeder_combout ),
	.Cout(),
	.Q(\macro_inst|serial_lim_input_inst|trigger_sync1~q ));
defparam \macro_inst|serial_lim_input_inst|trigger_sync1 .coord_x = 4;
defparam \macro_inst|serial_lim_input_inst|trigger_sync1 .coord_y = 4;
defparam \macro_inst|serial_lim_input_inst|trigger_sync1 .coord_z = 15;
defparam \macro_inst|serial_lim_input_inst|trigger_sync1 .mask = 16'hFF00;
defparam \macro_inst|serial_lim_input_inst|trigger_sync1 .modeMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|trigger_sync1 .FeedbackMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|trigger_sync1 .ShiftMux = 1'b0;
defparam \macro_inst|serial_lim_input_inst|trigger_sync1 .BypassEn = 1'b0;
defparam \macro_inst|serial_lim_input_inst|trigger_sync1 .CarryEnb = 1'b1;

alta_pllve \pll_inst|auto_generated|pll1 (
	.clkin(\PIN_HSE~input_o ),
	.clkfb(\pll_inst|auto_generated|pll1~FBOUT ),
	.pfden(vcc),
	.resetn(!\PLL_ENABLE~combout ),
	.phasecounterselect({gnd, gnd, gnd}),
	.phaseupdown(gnd),
	.phasestep(gnd),
	.scanclk(gnd),
	.scanclkena(vcc),
	.scandata(gnd),
	.configupdate(gnd),
	.scandataout(),
	.scandone(),
	.phasedone(),
	.clkout0(\pll_inst|auto_generated|pll1_CLK_bus [0]),
	.clkout1(\pll_inst|auto_generated|pll1_CLK_bus [1]),
	.clkout2(\pll_inst|auto_generated|pll1_CLK_bus [2]),
	.clkout3(\pll_inst|auto_generated|pll1_CLK_bus [3]),
	.clkout4(\pll_inst|auto_generated|pll1_CLK_bus [4]),
	.clkfbout(\pll_inst|auto_generated|pll1~FBOUT ),
	.lock(\auto_generated_inst.hbo_13_1bc039b416d3bc4a_bp ));
defparam \pll_inst|auto_generated|pll1 .coord_x = 22;
defparam \pll_inst|auto_generated|pll1 .coord_y = 5;
defparam \pll_inst|auto_generated|pll1 .coord_z = 0;
defparam \pll_inst|auto_generated|pll1 .CLKIN_HIGH = 8'b11111111;
defparam \pll_inst|auto_generated|pll1 .CLKIN_LOW = 8'b11111111;
defparam \pll_inst|auto_generated|pll1 .CLKIN_TRIM = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKIN_BYPASS = 1'b1;
defparam \pll_inst|auto_generated|pll1 .CLKFB_HIGH = 8'b00011101;
defparam \pll_inst|auto_generated|pll1 .CLKFB_LOW = 8'b00011101;
defparam \pll_inst|auto_generated|pll1 .CLKFB_TRIM = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKFB_BYPASS = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKDIV0_EN = 1'b1;
defparam \pll_inst|auto_generated|pll1 .CLKDIV1_EN = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKDIV2_EN = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKDIV3_EN = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKDIV4_EN = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT0_HIGH = 8'b00000010;
defparam \pll_inst|auto_generated|pll1 .CLKOUT0_LOW = 8'b00000010;
defparam \pll_inst|auto_generated|pll1 .CLKOUT0_TRIM = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT0_BYPASS = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT1_HIGH = 8'b11111111;
defparam \pll_inst|auto_generated|pll1 .CLKOUT1_LOW = 8'b11111111;
defparam \pll_inst|auto_generated|pll1 .CLKOUT1_TRIM = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT1_BYPASS = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT2_HIGH = 8'b11111111;
defparam \pll_inst|auto_generated|pll1 .CLKOUT2_LOW = 8'b11111111;
defparam \pll_inst|auto_generated|pll1 .CLKOUT2_TRIM = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT2_BYPASS = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT3_HIGH = 8'b11111111;
defparam \pll_inst|auto_generated|pll1 .CLKOUT3_LOW = 8'b11111111;
defparam \pll_inst|auto_generated|pll1 .CLKOUT3_TRIM = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT3_BYPASS = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT4_HIGH = 8'b11111111;
defparam \pll_inst|auto_generated|pll1 .CLKOUT4_LOW = 8'b11111111;
defparam \pll_inst|auto_generated|pll1 .CLKOUT4_TRIM = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT4_BYPASS = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT0_DEL = 8'b00000000;
defparam \pll_inst|auto_generated|pll1 .CLKOUT1_DEL = 8'b00000000;
defparam \pll_inst|auto_generated|pll1 .CLKOUT2_DEL = 8'b00000000;
defparam \pll_inst|auto_generated|pll1 .CLKOUT3_DEL = 8'b00000000;
defparam \pll_inst|auto_generated|pll1 .CLKOUT4_DEL = 8'b00000000;
defparam \pll_inst|auto_generated|pll1 .CLKOUT0_PHASE = 3'b000;
defparam \pll_inst|auto_generated|pll1 .CLKOUT1_PHASE = 3'b000;
defparam \pll_inst|auto_generated|pll1 .CLKOUT2_PHASE = 3'b000;
defparam \pll_inst|auto_generated|pll1 .CLKOUT3_PHASE = 3'b000;
defparam \pll_inst|auto_generated|pll1 .CLKOUT4_PHASE = 3'b000;
defparam \pll_inst|auto_generated|pll1 .CLKFB_DEL = 8'b00000000;
defparam \pll_inst|auto_generated|pll1 .CLKFB_PHASE = 3'b000;
defparam \pll_inst|auto_generated|pll1 .FEEDBACK_MODE = 3'b100;
defparam \pll_inst|auto_generated|pll1 .FBDELAY_VAL = 3'b100;
defparam \pll_inst|auto_generated|pll1 .PLLOUTP_EN = 1'b0;
defparam \pll_inst|auto_generated|pll1 .PLLOUTN_EN = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT1_CASCADE = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT2_CASCADE = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT3_CASCADE = 1'b0;
defparam \pll_inst|auto_generated|pll1 .CLKOUT4_CASCADE = 1'b0;
defparam \pll_inst|auto_generated|pll1 .VCO_POST_DIV = 1'b1;
defparam \pll_inst|auto_generated|pll1 .REG_CTRL = 2'b00;
defparam \pll_inst|auto_generated|pll1 .CP = 3'b100;
defparam \pll_inst|auto_generated|pll1 .RREF = 2'b01;
defparam \pll_inst|auto_generated|pll1 .RVI = 2'b01;
defparam \pll_inst|auto_generated|pll1 .IVCO = 3'b010;
defparam \pll_inst|auto_generated|pll1 .PLL_EN_FLAG = 1'b1;

alta_slice \pll_inst|auto_generated|pll_lock_sync (
	.A(vcc),
	.B(vcc),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(\pll_inst|auto_generated|pll_lock_sync~q ),
	.Clk(\auto_generated_inst.hbo_13_1bc039b416d3bc4a_bp_X48_Y1_SIG_VCC ),
	.AsyncReset(\PLL_ENABLE~clkctrl_outclk__AsyncReset_X48_Y1_SIG ),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\pll_inst|auto_generated|pll_lock_sync~feeder_combout ),
	.Cout(),
	.Q(\pll_inst|auto_generated|pll_lock_sync~q ));
defparam \pll_inst|auto_generated|pll_lock_sync .coord_x = 5;
defparam \pll_inst|auto_generated|pll_lock_sync .coord_y = 3;
defparam \pll_inst|auto_generated|pll_lock_sync .coord_z = 3;
defparam \pll_inst|auto_generated|pll_lock_sync .mask = 16'hFFFF;
defparam \pll_inst|auto_generated|pll_lock_sync .modeMux = 1'b0;
defparam \pll_inst|auto_generated|pll_lock_sync .FeedbackMux = 1'b0;
defparam \pll_inst|auto_generated|pll_lock_sync .ShiftMux = 1'b0;
defparam \pll_inst|auto_generated|pll_lock_sync .BypassEn = 1'b0;
defparam \pll_inst|auto_generated|pll_lock_sync .CarryEnb = 1'b1;

alta_rv32 rv32(
	.sys_clk(\gclksw_inst|gclk_switch__alta_gclksw__clkout ),
	.mem_ahb_hready(\rv32.mem_ahb_hready ),
	.mem_ahb_hreadyout(vcc),
	.mem_ahb_htrans({\rv32.mem_ahb_htrans[1] , \rv32.mem_ahb_htrans[0] }),
	.mem_ahb_hsize({\rv32.mem_ahb_hsize[2] , \rv32.mem_ahb_hsize[1] , \rv32.mem_ahb_hsize[0] }),
	.mem_ahb_hburst({\rv32.mem_ahb_hburst[2] , \rv32.mem_ahb_hburst[1] , \rv32.mem_ahb_hburst[0] }),
	.mem_ahb_hwrite(\rv32.mem_ahb_hwrite ),
	.mem_ahb_haddr({\rv32.mem_ahb_haddr[31] , \rv32.mem_ahb_haddr[30] , \rv32.mem_ahb_haddr[29] , \rv32.mem_ahb_haddr[28] , \rv32.mem_ahb_haddr[27] , \rv32.mem_ahb_haddr[26] , \rv32.mem_ahb_haddr[25] , \rv32.mem_ahb_haddr[24] , \rv32.mem_ahb_haddr[23] , \rv32.mem_ahb_haddr[22] , \rv32.mem_ahb_haddr[21] , \rv32.mem_ahb_haddr[20] , \rv32.mem_ahb_haddr[19] , \rv32.mem_ahb_haddr[18] , \rv32.mem_ahb_haddr[17] , \rv32.mem_ahb_haddr[16] , \rv32.mem_ahb_haddr[15] , \rv32.mem_ahb_haddr[14] , \rv32.mem_ahb_haddr[13] , \rv32.mem_ahb_haddr[12] , \rv32.mem_ahb_haddr[11] , \rv32.mem_ahb_haddr[10] , \rv32.mem_ahb_haddr[9] , \rv32.mem_ahb_haddr[8] , \rv32.mem_ahb_haddr[7] , \rv32.mem_ahb_haddr[6] , \rv32.mem_ahb_haddr[5] , \rv32.mem_ahb_haddr[4] , \rv32.mem_ahb_haddr[3] , \rv32.mem_ahb_haddr[2] , \rv32.mem_ahb_haddr[1] , \rv32.mem_ahb_haddr[0] }),
	.mem_ahb_hwdata({\rv32.mem_ahb_hwdata[31] , \rv32.mem_ahb_hwdata[30] , \rv32.mem_ahb_hwdata[29] , \rv32.mem_ahb_hwdata[28] , \rv32.mem_ahb_hwdata[27] , \rv32.mem_ahb_hwdata[26] , \rv32.mem_ahb_hwdata[25] , \rv32.mem_ahb_hwdata[24] , \rv32.mem_ahb_hwdata[23] , \rv32.mem_ahb_hwdata[22] , \rv32.mem_ahb_hwdata[21] , \rv32.mem_ahb_hwdata[20] , \rv32.mem_ahb_hwdata[19] , \rv32.mem_ahb_hwdata[18] , \rv32.mem_ahb_hwdata[17] , \rv32.mem_ahb_hwdata[16] , \rv32.mem_ahb_hwdata[15] , \rv32.mem_ahb_hwdata[14] , \rv32.mem_ahb_hwdata[13] , \rv32.mem_ahb_hwdata[12] , \rv32.mem_ahb_hwdata[11] , \rv32.mem_ahb_hwdata[10] , \rv32.mem_ahb_hwdata[9] , \rv32.mem_ahb_hwdata[8] , \rv32.mem_ahb_hwdata[7] , \rv32.mem_ahb_hwdata[6] , \rv32.mem_ahb_hwdata[5] , \rv32.mem_ahb_hwdata[4] , \rv32.mem_ahb_hwdata[3] , \rv32.mem_ahb_hwdata[2] , \rv32.mem_ahb_hwdata[1] , \rv32.mem_ahb_hwdata[0] }),
	.mem_ahb_hresp(gnd),
	.mem_ahb_hrdata({\macro_inst|mem_ahb_hrdata[31]~31_combout , \macro_inst|mem_ahb_hrdata[30]~30_combout , \macro_inst|mem_ahb_hrdata[29]~29_combout , \macro_inst|mem_ahb_hrdata[28]~28_combout , \macro_inst|mem_ahb_hrdata[27]~27_combout , \macro_inst|mem_ahb_hrdata[26]~26_combout , \macro_inst|mem_ahb_hrdata[25]~25_combout , \macro_inst|mem_ahb_hrdata[24]~24_combout , \macro_inst|mem_ahb_hrdata[23]~23_combout , \macro_inst|mem_ahb_hrdata[22]~22_combout , \macro_inst|mem_ahb_hrdata[21]~21_combout , \macro_inst|mem_ahb_hrdata[20]~20_combout , \macro_inst|mem_ahb_hrdata[19]~19_combout , \macro_inst|mem_ahb_hrdata[18]~18_combout , \macro_inst|mem_ahb_hrdata[17]~17_combout , \macro_inst|mem_ahb_hrdata[16]~16_combout , \macro_inst|mem_ahb_hrdata[15]~15_combout , \macro_inst|mem_ahb_hrdata[14]~14_combout , \macro_inst|mem_ahb_hrdata[13]~13_combout , \macro_inst|mem_ahb_hrdata[12]~12_combout , \macro_inst|mem_ahb_hrdata[11]~11_combout , \macro_inst|mem_ahb_hrdata[10]~10_combout , \macro_inst|mem_ahb_hrdata[9]~9_combout , \macro_inst|mem_ahb_hrdata[8]~8_combout , \macro_inst|mem_ahb_hrdata[7]~7_combout , \macro_inst|mem_ahb_hrdata[6]~6_combout , \macro_inst|mem_ahb_hrdata[5]~5_combout , \macro_inst|mem_ahb_hrdata[4]~4_combout , \macro_inst|mem_ahb_hrdata[3]~3_combout , \macro_inst|mem_ahb_hrdata[2]~2_combout , \macro_inst|mem_ahb_hrdata[1]~1_combout , \macro_inst|mem_ahb_hrdata[0]~0_combout }),
	.slave_ahb_hsel(gnd),
	.slave_ahb_hready(vcc),
	.slave_ahb_hreadyout(\rv32.slave_ahb_hreadyout ),
	.slave_ahb_htrans({gnd, gnd}),
	.slave_ahb_hsize({gnd, gnd, gnd}),
	.slave_ahb_hburst({gnd, gnd, gnd}),
	.slave_ahb_hwrite(gnd),
	.slave_ahb_haddr({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
	.slave_ahb_hwdata({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
	.slave_ahb_hresp(\rv32.slave_ahb_hresp ),
	.slave_ahb_hrdata({\rv32.slave_ahb_hrdata[31] , \rv32.slave_ahb_hrdata[30] , \rv32.slave_ahb_hrdata[29] , \rv32.slave_ahb_hrdata[28] , \rv32.slave_ahb_hrdata[27] , \rv32.slave_ahb_hrdata[26] , \rv32.slave_ahb_hrdata[25] , \rv32.slave_ahb_hrdata[24] , \rv32.slave_ahb_hrdata[23] , \rv32.slave_ahb_hrdata[22] , \rv32.slave_ahb_hrdata[21] , \rv32.slave_ahb_hrdata[20] , \rv32.slave_ahb_hrdata[19] , \rv32.slave_ahb_hrdata[18] , \rv32.slave_ahb_hrdata[17] , \rv32.slave_ahb_hrdata[16] , \rv32.slave_ahb_hrdata[15] , \rv32.slave_ahb_hrdata[14] , \rv32.slave_ahb_hrdata[13] , \rv32.slave_ahb_hrdata[12] , \rv32.slave_ahb_hrdata[11] , \rv32.slave_ahb_hrdata[10] , \rv32.slave_ahb_hrdata[9] , \rv32.slave_ahb_hrdata[8] , \rv32.slave_ahb_hrdata[7] , \rv32.slave_ahb_hrdata[6] , \rv32.slave_ahb_hrdata[5] , \rv32.slave_ahb_hrdata[4] , \rv32.slave_ahb_hrdata[3] , \rv32.slave_ahb_hrdata[2] , \rv32.slave_ahb_hrdata[1] , \rv32.slave_ahb_hrdata[0] }),
	.gpio0_io_in({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
	.gpio0_io_out_data({\rv32.gpio0_io_out_data[7] , \rv32.gpio0_io_out_data[6] , \rv32.gpio0_io_out_data[5] , \rv32.gpio0_io_out_data[4] , \rv32.gpio0_io_out_data[3] , \rv32.gpio0_io_out_data[2] , \rv32.gpio0_io_out_data[1] , \rv32.gpio0_io_out_data[0] }),
	.gpio0_io_out_en({\rv32.gpio0_io_out_en[7] , \rv32.gpio0_io_out_en[6] , \rv32.gpio0_io_out_en[5] , \rv32.gpio0_io_out_en[4] , \rv32.gpio0_io_out_en[3] , \rv32.gpio0_io_out_en[2] , \rv32.gpio0_io_out_en[1] , \rv32.gpio0_io_out_en[0] }),
	.gpio1_io_in({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
	.gpio1_io_out_data({\rv32.gpio1_io_out_data[7] , \rv32.gpio1_io_out_data[6] , \rv32.gpio1_io_out_data[5] , \rv32.gpio1_io_out_data[4] , \rv32.gpio1_io_out_data[3] , \rv32.gpio1_io_out_data[2] , \rv32.gpio1_io_out_data[1] , \rv32.gpio1_io_out_data[0] }),
	.gpio1_io_out_en({\rv32.gpio1_io_out_en[7] , \rv32.gpio1_io_out_en[6] , \rv32.gpio1_io_out_en[5] , \rv32.gpio1_io_out_en[4] , \rv32.gpio1_io_out_en[3] , \rv32.gpio1_io_out_en[2] , \rv32.gpio1_io_out_en[1] , \rv32.gpio1_io_out_en[0] }),
	.sys_ctrl_clkSource({\rv32.sys_ctrl_clkSource[1] , \rv32.sys_ctrl_clkSource[0] }),
	.sys_ctrl_hseEnable(\rv32.sys_ctrl_hseEnable ),
	.sys_ctrl_hseBypass(\rv32.sys_ctrl_hseBypass ),
	.sys_ctrl_pllEnable(\rv32.sys_ctrl_pllEnable ),
	.sys_ctrl_pllReady(\auto_generated_inst.hbo_13_1bc039b416d3bc4a_bp ),
	.sys_ctrl_sleep(\rv32.sys_ctrl_sleep ),
	.sys_ctrl_stop(\rv32.sys_ctrl_stop ),
	.sys_ctrl_standby(\rv32.sys_ctrl_standby ),
	.gpio2_io_in({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
	.gpio2_io_out_data({\rv32.gpio2_io_out_data[7] , \rv32.gpio2_io_out_data[6] , \rv32.gpio2_io_out_data[5] , \rv32.gpio2_io_out_data[4] , \rv32.gpio2_io_out_data[3] , \rv32.gpio2_io_out_data[2] , \rv32.gpio2_io_out_data[1] , \rv32.gpio2_io_out_data[0] }),
	.gpio2_io_out_en({\rv32.gpio2_io_out_en[7] , \rv32.gpio2_io_out_en[6] , \rv32.gpio2_io_out_en[5] , \rv32.gpio2_io_out_en[4] , \rv32.gpio2_io_out_en[3] , \rv32.gpio2_io_out_en[2] , \rv32.gpio2_io_out_en[1] , \rv32.gpio2_io_out_en[0] }),
	.gpio3_io_in({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
	.gpio3_io_out_data({\rv32.gpio3_io_out_data[7] , \rv32.gpio3_io_out_data[6] , \rv32.gpio3_io_out_data[5] , \rv32.gpio3_io_out_data[4] , \rv32.gpio3_io_out_data[3] , \rv32.gpio3_io_out_data[2] , \rv32.gpio3_io_out_data[1] , \rv32.gpio3_io_out_data[0] }),
	.gpio3_io_out_en({\rv32.gpio3_io_out_en[7] , \rv32.gpio3_io_out_en[6] , \rv32.gpio3_io_out_en[5] , \rv32.gpio3_io_out_en[4] , \rv32.gpio3_io_out_en[3] , \rv32.gpio3_io_out_en[2] , \rv32.gpio3_io_out_en[1] , \rv32.gpio3_io_out_en[0] }),
	.gpio4_io_in({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
	.gpio4_io_out_data({\rv32.gpio4_io_out_data[7] , \rv32.gpio4_io_out_data[6] , \rv32.gpio4_io_out_data[5] , \rv32.gpio4_io_out_data[4] , \rv32.gpio4_io_out_data[3] , \rv32.gpio4_io_out_data[2] , \rv32.gpio4_io_out_data[1] , \rv32.gpio4_io_out_data[0] }),
	.gpio4_io_out_en({\rv32.gpio4_io_out_en[7] , \rv32.gpio4_io_out_en[6] , \rv32.gpio4_io_out_en[5] , \rv32.gpio4_io_out_en[4] , \rv32.gpio4_io_out_en[3] , \rv32.gpio4_io_out_en[2] , \rv32.gpio4_io_out_en[1] , \rv32.gpio4_io_out_en[0] }),
	.gpio5_io_in({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
	.gpio5_io_out_data({\rv32.gpio5_io_out_data[7] , \rv32.gpio5_io_out_data[6] , \rv32.gpio5_io_out_data[5] , \rv32.gpio5_io_out_data[4] , \rv32.gpio5_io_out_data[3] , \rv32.gpio5_io_out_data[2] , \rv32.gpio5_io_out_data[1] , \rv32.gpio5_io_out_data[0] }),
	.gpio5_io_out_en({\rv32.gpio5_io_out_en[7] , \rv32.gpio5_io_out_en[6] , \rv32.gpio5_io_out_en[5] , \rv32.gpio5_io_out_en[4] , \rv32.gpio5_io_out_en[3] , \rv32.gpio5_io_out_en[2] , \rv32.gpio5_io_out_en[1] , \rv32.gpio5_io_out_en[0] }),
	.gpio6_io_in({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
	.gpio6_io_out_data({\rv32.gpio6_io_out_data[7] , \rv32.gpio6_io_out_data[6] , \rv32.gpio6_io_out_data[5] , \rv32.gpio6_io_out_data[4] , \rv32.gpio6_io_out_data[3] , \rv32.gpio6_io_out_data[2] , \rv32.gpio6_io_out_data[1] , \rv32.gpio6_io_out_data[0] }),
	.gpio6_io_out_en({\rv32.gpio6_io_out_en[7] , \rv32.gpio6_io_out_en[6] , \rv32.gpio6_io_out_en[5] , \rv32.gpio6_io_out_en[4] , \rv32.gpio6_io_out_en[3] , \rv32.gpio6_io_out_en[2] , \rv32.gpio6_io_out_en[1] , \rv32.gpio6_io_out_en[0] }),
	.gpio7_io_in({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
	.gpio7_io_out_data({\rv32.gpio7_io_out_data[7] , \rv32.gpio7_io_out_data[6] , \rv32.gpio7_io_out_data[5] , \rv32.gpio7_io_out_data[4] , \rv32.gpio7_io_out_data[3] , \rv32.gpio7_io_out_data[2] , \rv32.gpio7_io_out_data[1] , \rv32.gpio7_io_out_data[0] }),
	.gpio7_io_out_en({\rv32.gpio7_io_out_en[7] , \rv32.gpio7_io_out_en[6] , \rv32.gpio7_io_out_en[5] , \rv32.gpio7_io_out_en[4] , \rv32.gpio7_io_out_en[3] , \rv32.gpio7_io_out_en[2] , \rv32.gpio7_io_out_en[1] , \rv32.gpio7_io_out_en[0] }),
	.gpio8_io_in({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
	.gpio8_io_out_data({\rv32.gpio8_io_out_data[7] , \rv32.gpio8_io_out_data[6] , \rv32.gpio8_io_out_data[5] , \rv32.gpio8_io_out_data[4] , \rv32.gpio8_io_out_data[3] , \rv32.gpio8_io_out_data[2] , \rv32.gpio8_io_out_data[1] , \rv32.gpio8_io_out_data[0] }),
	.gpio8_io_out_en({\rv32.gpio8_io_out_en[7] , \rv32.gpio8_io_out_en[6] , \rv32.gpio8_io_out_en[5] , \rv32.gpio8_io_out_en[4] , \rv32.gpio8_io_out_en[3] , \rv32.gpio8_io_out_en[2] , \rv32.gpio8_io_out_en[1] , \rv32.gpio8_io_out_en[0] }),
	.gpio9_io_in({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
	.gpio9_io_out_data({\rv32.gpio9_io_out_data[7] , \rv32.gpio9_io_out_data[6] , \rv32.gpio9_io_out_data[5] , \rv32.gpio9_io_out_data[4] , \rv32.gpio9_io_out_data[3] , \rv32.gpio9_io_out_data[2] , \rv32.gpio9_io_out_data[1] , \rv32.gpio9_io_out_data[0] }),
	.gpio9_io_out_en({\rv32.gpio9_io_out_en[7] , \rv32.gpio9_io_out_en[6] , \rv32.gpio9_io_out_en[5] , \rv32.gpio9_io_out_en[4] , \rv32.gpio9_io_out_en[3] , \rv32.gpio9_io_out_en[2] , \rv32.gpio9_io_out_en[1] , \rv32.gpio9_io_out_en[0] }),
	.ext_resetn(vcc),
	.resetn_out(\rv32.resetn_out ),
	.dmactive(\rv32.dmactive ),
	.swj_JTAGNSW(\rv32.swj_JTAGNSW ),
	.swj_JTAGSTATE({\rv32.swj_JTAGSTATE[3] , \rv32.swj_JTAGSTATE[2] , \rv32.swj_JTAGSTATE[1] , \rv32.swj_JTAGSTATE[0] }),
	.swj_JTAGIR({\rv32.swj_JTAGIR[3] , \rv32.swj_JTAGIR[2] , \rv32.swj_JTAGIR[1] , \rv32.swj_JTAGIR[0] }),
	.ext_int({gnd, gnd, gnd, gnd, gnd, gnd, gnd, gnd}),
	.ext_dma_DMACBREQ({gnd, gnd, gnd, gnd}),
	.ext_dma_DMACLBREQ({gnd, gnd, gnd, gnd}),
	.ext_dma_DMACSREQ({gnd, gnd, gnd, gnd}),
	.ext_dma_DMACLSREQ({gnd, gnd, gnd, gnd}),
	.ext_dma_DMACCLR({\rv32.ext_dma_DMACCLR[3] , \rv32.ext_dma_DMACCLR[2] , \rv32.ext_dma_DMACCLR[1] , \rv32.ext_dma_DMACCLR[0] }),
	.ext_dma_DMACTC({\rv32.ext_dma_DMACTC[3] , \rv32.ext_dma_DMACTC[2] , \rv32.ext_dma_DMACTC[1] , \rv32.ext_dma_DMACTC[0] }),
	.local_int({gnd, gnd, gnd, gnd}),
	.test_mode({gnd, gnd}),
	.usb0_xcvr_clk(vcc),
	.usb0_id(vcc));
defparam rv32.coord_x = 0;
defparam rv32.coord_y = 5;
defparam rv32.coord_z = 0;

alta_syncctrl syncload_ctrl_X43_Y2(
	.Din(),
	.Dout(SyncLoad_X43_Y2_GND));
defparam syncload_ctrl_X43_Y2.coord_x = 7;
defparam syncload_ctrl_X43_Y2.coord_y = 2;
defparam syncload_ctrl_X43_Y2.coord_z = 1;
defparam syncload_ctrl_X43_Y2.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X46_Y2(
	.Din(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q ),
	.Dout(\macro_inst|serial_lim_input_inst|state_reg.STATE_LOAD~q__SyncLoad_X46_Y2_INV ));
defparam syncload_ctrl_X46_Y2.coord_x = 4;
defparam syncload_ctrl_X46_Y2.coord_y = 3;
defparam syncload_ctrl_X46_Y2.coord_z = 1;
defparam syncload_ctrl_X46_Y2.SyncCtrlMux = 2'b11;

alta_syncctrl syncload_ctrl_X46_Y3(
	.Din(),
	.Dout(SyncLoad_X46_Y3_VCC));
defparam syncload_ctrl_X46_Y3.coord_x = 5;
defparam syncload_ctrl_X46_Y3.coord_y = 4;
defparam syncload_ctrl_X46_Y3.coord_z = 1;
defparam syncload_ctrl_X46_Y3.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X47_Y3(
	.Din(),
	.Dout(SyncLoad_X47_Y3_VCC));
defparam syncload_ctrl_X47_Y3.coord_x = 4;
defparam syncload_ctrl_X47_Y3.coord_y = 4;
defparam syncload_ctrl_X47_Y3.coord_z = 1;
defparam syncload_ctrl_X47_Y3.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X49_Y2(
	.Din(),
	.Dout(SyncLoad_X49_Y2_VCC));
defparam syncload_ctrl_X49_Y2.coord_x = 9;
defparam syncload_ctrl_X49_Y2.coord_y = 3;
defparam syncload_ctrl_X49_Y2.coord_z = 1;
defparam syncload_ctrl_X49_Y2.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X49_Y3(
	.Din(),
	.Dout(SyncLoad_X49_Y3_VCC));
defparam syncload_ctrl_X49_Y3.coord_x = 6;
defparam syncload_ctrl_X49_Y3.coord_y = 4;
defparam syncload_ctrl_X49_Y3.coord_z = 1;
defparam syncload_ctrl_X49_Y3.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X50_Y1(
	.Din(\macro_inst|controller|serial|state.IDLE~q ),
	.Dout(\macro_inst|controller|serial|state.IDLE~q__SyncLoad_X50_Y1_INV ));
defparam syncload_ctrl_X50_Y1.coord_x = 7;
defparam syncload_ctrl_X50_Y1.coord_y = 1;
defparam syncload_ctrl_X50_Y1.coord_z = 1;
defparam syncload_ctrl_X50_Y1.SyncCtrlMux = 2'b11;

alta_syncctrl syncload_ctrl_X50_Y2(
	.Din(),
	.Dout(SyncLoad_X50_Y2_GND));
defparam syncload_ctrl_X50_Y2.coord_x = 9;
defparam syncload_ctrl_X50_Y2.coord_y = 2;
defparam syncload_ctrl_X50_Y2.coord_z = 1;
defparam syncload_ctrl_X50_Y2.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X50_Y3(
	.Din(),
	.Dout(SyncLoad_X50_Y3_VCC));
defparam syncload_ctrl_X50_Y3.coord_x = 8;
defparam syncload_ctrl_X50_Y3.coord_y = 4;
defparam syncload_ctrl_X50_Y3.coord_z = 1;
defparam syncload_ctrl_X50_Y3.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X51_Y2(
	.Din(),
	.Dout(SyncLoad_X51_Y2_GND));
defparam syncload_ctrl_X51_Y2.coord_x = 8;
defparam syncload_ctrl_X51_Y2.coord_y = 2;
defparam syncload_ctrl_X51_Y2.coord_z = 1;
defparam syncload_ctrl_X51_Y2.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X51_Y3(
	.Din(),
	.Dout(SyncLoad_X51_Y3_VCC));
defparam syncload_ctrl_X51_Y3.coord_x = 9;
defparam syncload_ctrl_X51_Y3.coord_y = 4;
defparam syncload_ctrl_X51_Y3.coord_z = 1;
defparam syncload_ctrl_X51_Y3.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X51_Y4(
	.Din(),
	.Dout(SyncLoad_X51_Y4_VCC));
defparam syncload_ctrl_X51_Y4.coord_x = 15;
defparam syncload_ctrl_X51_Y4.coord_y = 2;
defparam syncload_ctrl_X51_Y4.coord_z = 1;
defparam syncload_ctrl_X51_Y4.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X52_Y2(
	.Din(),
	.Dout(SyncLoad_X52_Y2_VCC));
defparam syncload_ctrl_X52_Y2.coord_x = 16;
defparam syncload_ctrl_X52_Y2.coord_y = 5;
defparam syncload_ctrl_X52_Y2.coord_z = 1;
defparam syncload_ctrl_X52_Y2.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X52_Y3(
	.Din(),
	.Dout(SyncLoad_X52_Y3_VCC));
defparam syncload_ctrl_X52_Y3.coord_x = 8;
defparam syncload_ctrl_X52_Y3.coord_y = 3;
defparam syncload_ctrl_X52_Y3.coord_z = 1;
defparam syncload_ctrl_X52_Y3.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X52_Y4(
	.Din(),
	.Dout(SyncLoad_X52_Y4_VCC));
defparam syncload_ctrl_X52_Y4.coord_x = 16;
defparam syncload_ctrl_X52_Y4.coord_y = 2;
defparam syncload_ctrl_X52_Y4.coord_z = 1;
defparam syncload_ctrl_X52_Y4.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X53_Y4(
	.Din(),
	.Dout(SyncLoad_X53_Y4_VCC));
defparam syncload_ctrl_X53_Y4.coord_x = 15;
defparam syncload_ctrl_X53_Y4.coord_y = 4;
defparam syncload_ctrl_X53_Y4.coord_z = 1;
defparam syncload_ctrl_X53_Y4.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X54_Y1(
	.Din(),
	.Dout(SyncLoad_X54_Y1_VCC));
defparam syncload_ctrl_X54_Y1.coord_x = 20;
defparam syncload_ctrl_X54_Y1.coord_y = 2;
defparam syncload_ctrl_X54_Y1.coord_z = 1;
defparam syncload_ctrl_X54_Y1.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X54_Y2(
	.Din(),
	.Dout(SyncLoad_X54_Y2_VCC));
defparam syncload_ctrl_X54_Y2.coord_x = 14;
defparam syncload_ctrl_X54_Y2.coord_y = 5;
defparam syncload_ctrl_X54_Y2.coord_z = 1;
defparam syncload_ctrl_X54_Y2.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X54_Y3(
	.Din(),
	.Dout(SyncLoad_X54_Y3_VCC));
defparam syncload_ctrl_X54_Y3.coord_x = 14;
defparam syncload_ctrl_X54_Y3.coord_y = 12;
defparam syncload_ctrl_X54_Y3.coord_z = 1;
defparam syncload_ctrl_X54_Y3.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X54_Y4(
	.Din(),
	.Dout(SyncLoad_X54_Y4_VCC));
defparam syncload_ctrl_X54_Y4.coord_x = 11;
defparam syncload_ctrl_X54_Y4.coord_y = 2;
defparam syncload_ctrl_X54_Y4.coord_z = 1;
defparam syncload_ctrl_X54_Y4.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X56_Y1(
	.Din(),
	.Dout(SyncLoad_X56_Y1_VCC));
defparam syncload_ctrl_X56_Y1.coord_x = 10;
defparam syncload_ctrl_X56_Y1.coord_y = 2;
defparam syncload_ctrl_X56_Y1.coord_z = 1;
defparam syncload_ctrl_X56_Y1.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X56_Y10(
	.Din(),
	.Dout(SyncLoad_X56_Y10_VCC));
defparam syncload_ctrl_X56_Y10.coord_x = 11;
defparam syncload_ctrl_X56_Y10.coord_y = 3;
defparam syncload_ctrl_X56_Y10.coord_z = 1;
defparam syncload_ctrl_X56_Y10.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X56_Y2(
	.Din(),
	.Dout(SyncLoad_X56_Y2_VCC));
defparam syncload_ctrl_X56_Y2.coord_x = 16;
defparam syncload_ctrl_X56_Y2.coord_y = 11;
defparam syncload_ctrl_X56_Y2.coord_z = 1;
defparam syncload_ctrl_X56_Y2.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X56_Y3(
	.Din(),
	.Dout(SyncLoad_X56_Y3_GND));
defparam syncload_ctrl_X56_Y3.coord_x = 12;
defparam syncload_ctrl_X56_Y3.coord_y = 4;
defparam syncload_ctrl_X56_Y3.coord_z = 1;
defparam syncload_ctrl_X56_Y3.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X56_Y4(
	.Din(),
	.Dout(SyncLoad_X56_Y4_VCC));
defparam syncload_ctrl_X56_Y4.coord_x = 17;
defparam syncload_ctrl_X56_Y4.coord_y = 4;
defparam syncload_ctrl_X56_Y4.coord_z = 1;
defparam syncload_ctrl_X56_Y4.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X56_Y5(
	.Din(),
	.Dout(SyncLoad_X56_Y5_GND));
defparam syncload_ctrl_X56_Y5.coord_x = 10;
defparam syncload_ctrl_X56_Y5.coord_y = 4;
defparam syncload_ctrl_X56_Y5.coord_z = 1;
defparam syncload_ctrl_X56_Y5.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X56_Y6(
	.Din(),
	.Dout(SyncLoad_X56_Y6_VCC));
defparam syncload_ctrl_X56_Y6.coord_x = 17;
defparam syncload_ctrl_X56_Y6.coord_y = 2;
defparam syncload_ctrl_X56_Y6.coord_z = 1;
defparam syncload_ctrl_X56_Y6.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X56_Y7(
	.Din(),
	.Dout(SyncLoad_X56_Y7_VCC));
defparam syncload_ctrl_X56_Y7.coord_x = 14;
defparam syncload_ctrl_X56_Y7.coord_y = 2;
defparam syncload_ctrl_X56_Y7.coord_z = 1;
defparam syncload_ctrl_X56_Y7.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X56_Y8(
	.Din(),
	.Dout(SyncLoad_X56_Y8_VCC));
defparam syncload_ctrl_X56_Y8.coord_x = 19;
defparam syncload_ctrl_X56_Y8.coord_y = 1;
defparam syncload_ctrl_X56_Y8.coord_z = 1;
defparam syncload_ctrl_X56_Y8.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X56_Y9(
	.Din(),
	.Dout(SyncLoad_X56_Y9_VCC));
defparam syncload_ctrl_X56_Y9.coord_x = 17;
defparam syncload_ctrl_X56_Y9.coord_y = 9;
defparam syncload_ctrl_X56_Y9.coord_z = 1;
defparam syncload_ctrl_X56_Y9.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X57_Y1(
	.Din(),
	.Dout(SyncLoad_X57_Y1_VCC));
defparam syncload_ctrl_X57_Y1.coord_x = 12;
defparam syncload_ctrl_X57_Y1.coord_y = 2;
defparam syncload_ctrl_X57_Y1.coord_z = 1;
defparam syncload_ctrl_X57_Y1.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X57_Y10(
	.Din(),
	.Dout(SyncLoad_X57_Y10_VCC));
defparam syncload_ctrl_X57_Y10.coord_x = 12;
defparam syncload_ctrl_X57_Y10.coord_y = 3;
defparam syncload_ctrl_X57_Y10.coord_z = 1;
defparam syncload_ctrl_X57_Y10.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X57_Y11(
	.Din(),
	.Dout(SyncLoad_X57_Y11_VCC));
defparam syncload_ctrl_X57_Y11.coord_x = 20;
defparam syncload_ctrl_X57_Y11.coord_y = 10;
defparam syncload_ctrl_X57_Y11.coord_z = 1;
defparam syncload_ctrl_X57_Y11.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X57_Y12(
	.Din(),
	.Dout(SyncLoad_X57_Y12_VCC));
defparam syncload_ctrl_X57_Y12.coord_x = 18;
defparam syncload_ctrl_X57_Y12.coord_y = 8;
defparam syncload_ctrl_X57_Y12.coord_z = 1;
defparam syncload_ctrl_X57_Y12.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X57_Y2(
	.Din(),
	.Dout(SyncLoad_X57_Y2_VCC));
defparam syncload_ctrl_X57_Y2.coord_x = 18;
defparam syncload_ctrl_X57_Y2.coord_y = 12;
defparam syncload_ctrl_X57_Y2.coord_z = 1;
defparam syncload_ctrl_X57_Y2.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X57_Y3(
	.Din(),
	.Dout(SyncLoad_X57_Y3_VCC));
defparam syncload_ctrl_X57_Y3.coord_x = 14;
defparam syncload_ctrl_X57_Y3.coord_y = 11;
defparam syncload_ctrl_X57_Y3.coord_z = 1;
defparam syncload_ctrl_X57_Y3.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X57_Y4(
	.Din(),
	.Dout(SyncLoad_X57_Y4_VCC));
defparam syncload_ctrl_X57_Y4.coord_x = 16;
defparam syncload_ctrl_X57_Y4.coord_y = 4;
defparam syncload_ctrl_X57_Y4.coord_z = 1;
defparam syncload_ctrl_X57_Y4.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X57_Y5(
	.Din(),
	.Dout(SyncLoad_X57_Y5_GND));
defparam syncload_ctrl_X57_Y5.coord_x = 14;
defparam syncload_ctrl_X57_Y5.coord_y = 7;
defparam syncload_ctrl_X57_Y5.coord_z = 1;
defparam syncload_ctrl_X57_Y5.SyncCtrlMux = 2'b00;

alta_syncctrl syncload_ctrl_X57_Y6(
	.Din(),
	.Dout(SyncLoad_X57_Y6_VCC));
defparam syncload_ctrl_X57_Y6.coord_x = 14;
defparam syncload_ctrl_X57_Y6.coord_y = 10;
defparam syncload_ctrl_X57_Y6.coord_z = 1;
defparam syncload_ctrl_X57_Y6.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X57_Y8(
	.Din(),
	.Dout(SyncLoad_X57_Y8_VCC));
defparam syncload_ctrl_X57_Y8.coord_x = 18;
defparam syncload_ctrl_X57_Y8.coord_y = 3;
defparam syncload_ctrl_X57_Y8.coord_z = 1;
defparam syncload_ctrl_X57_Y8.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X57_Y9(
	.Din(),
	.Dout(SyncLoad_X57_Y9_VCC));
defparam syncload_ctrl_X57_Y9.coord_x = 16;
defparam syncload_ctrl_X57_Y9.coord_y = 9;
defparam syncload_ctrl_X57_Y9.coord_z = 1;
defparam syncload_ctrl_X57_Y9.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X58_Y1(
	.Din(),
	.Dout(SyncLoad_X58_Y1_VCC));
defparam syncload_ctrl_X58_Y1.coord_x = 10;
defparam syncload_ctrl_X58_Y1.coord_y = 1;
defparam syncload_ctrl_X58_Y1.coord_z = 1;
defparam syncload_ctrl_X58_Y1.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X58_Y10(
	.Din(),
	.Dout(SyncLoad_X58_Y10_VCC));
defparam syncload_ctrl_X58_Y10.coord_x = 17;
defparam syncload_ctrl_X58_Y10.coord_y = 7;
defparam syncload_ctrl_X58_Y10.coord_z = 1;
defparam syncload_ctrl_X58_Y10.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X58_Y11(
	.Din(),
	.Dout(SyncLoad_X58_Y11_VCC));
defparam syncload_ctrl_X58_Y11.coord_x = 19;
defparam syncload_ctrl_X58_Y11.coord_y = 12;
defparam syncload_ctrl_X58_Y11.coord_z = 1;
defparam syncload_ctrl_X58_Y11.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X58_Y12(
	.Din(),
	.Dout(SyncLoad_X58_Y12_VCC));
defparam syncload_ctrl_X58_Y12.coord_x = 20;
defparam syncload_ctrl_X58_Y12.coord_y = 3;
defparam syncload_ctrl_X58_Y12.coord_z = 1;
defparam syncload_ctrl_X58_Y12.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X58_Y2(
	.Din(),
	.Dout(SyncLoad_X58_Y2_VCC));
defparam syncload_ctrl_X58_Y2.coord_x = 16;
defparam syncload_ctrl_X58_Y2.coord_y = 10;
defparam syncload_ctrl_X58_Y2.coord_z = 1;
defparam syncload_ctrl_X58_Y2.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X58_Y3(
	.Din(),
	.Dout(SyncLoad_X58_Y3_VCC));
defparam syncload_ctrl_X58_Y3.coord_x = 15;
defparam syncload_ctrl_X58_Y3.coord_y = 11;
defparam syncload_ctrl_X58_Y3.coord_z = 1;
defparam syncload_ctrl_X58_Y3.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X58_Y4(
	.Din(),
	.Dout(SyncLoad_X58_Y4_VCC));
defparam syncload_ctrl_X58_Y4.coord_x = 16;
defparam syncload_ctrl_X58_Y4.coord_y = 8;
defparam syncload_ctrl_X58_Y4.coord_z = 1;
defparam syncload_ctrl_X58_Y4.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X58_Y5(
	.Din(),
	.Dout(SyncLoad_X58_Y5_VCC));
defparam syncload_ctrl_X58_Y5.coord_x = 16;
defparam syncload_ctrl_X58_Y5.coord_y = 12;
defparam syncload_ctrl_X58_Y5.coord_z = 1;
defparam syncload_ctrl_X58_Y5.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X58_Y6(
	.Din(),
	.Dout(SyncLoad_X58_Y6_VCC));
defparam syncload_ctrl_X58_Y6.coord_x = 14;
defparam syncload_ctrl_X58_Y6.coord_y = 9;
defparam syncload_ctrl_X58_Y6.coord_z = 1;
defparam syncload_ctrl_X58_Y6.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X58_Y7(
	.Din(),
	.Dout(SyncLoad_X58_Y7_VCC));
defparam syncload_ctrl_X58_Y7.coord_x = 14;
defparam syncload_ctrl_X58_Y7.coord_y = 4;
defparam syncload_ctrl_X58_Y7.coord_z = 1;
defparam syncload_ctrl_X58_Y7.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X58_Y8(
	.Din(),
	.Dout(SyncLoad_X58_Y8_VCC));
defparam syncload_ctrl_X58_Y8.coord_x = 17;
defparam syncload_ctrl_X58_Y8.coord_y = 5;
defparam syncload_ctrl_X58_Y8.coord_z = 1;
defparam syncload_ctrl_X58_Y8.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X58_Y9(
	.Din(),
	.Dout(SyncLoad_X58_Y9_VCC));
defparam syncload_ctrl_X58_Y9.coord_x = 18;
defparam syncload_ctrl_X58_Y9.coord_y = 9;
defparam syncload_ctrl_X58_Y9.coord_z = 1;
defparam syncload_ctrl_X58_Y9.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X59_Y1(
	.Din(),
	.Dout(SyncLoad_X59_Y1_VCC));
defparam syncload_ctrl_X59_Y1.coord_x = 16;
defparam syncload_ctrl_X59_Y1.coord_y = 3;
defparam syncload_ctrl_X59_Y1.coord_z = 1;
defparam syncload_ctrl_X59_Y1.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X59_Y10(
	.Din(),
	.Dout(SyncLoad_X59_Y10_VCC));
defparam syncload_ctrl_X59_Y10.coord_x = 18;
defparam syncload_ctrl_X59_Y10.coord_y = 6;
defparam syncload_ctrl_X59_Y10.coord_z = 1;
defparam syncload_ctrl_X59_Y10.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X59_Y11(
	.Din(),
	.Dout(SyncLoad_X59_Y11_VCC));
defparam syncload_ctrl_X59_Y11.coord_x = 19;
defparam syncload_ctrl_X59_Y11.coord_y = 3;
defparam syncload_ctrl_X59_Y11.coord_z = 1;
defparam syncload_ctrl_X59_Y11.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X59_Y12(
	.Din(),
	.Dout(SyncLoad_X59_Y12_VCC));
defparam syncload_ctrl_X59_Y12.coord_x = 20;
defparam syncload_ctrl_X59_Y12.coord_y = 5;
defparam syncload_ctrl_X59_Y12.coord_z = 1;
defparam syncload_ctrl_X59_Y12.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X59_Y2(
	.Din(),
	.Dout(SyncLoad_X59_Y2_VCC));
defparam syncload_ctrl_X59_Y2.coord_x = 10;
defparam syncload_ctrl_X59_Y2.coord_y = 3;
defparam syncload_ctrl_X59_Y2.coord_z = 1;
defparam syncload_ctrl_X59_Y2.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X59_Y3(
	.Din(),
	.Dout(SyncLoad_X59_Y3_VCC));
defparam syncload_ctrl_X59_Y3.coord_x = 15;
defparam syncload_ctrl_X59_Y3.coord_y = 12;
defparam syncload_ctrl_X59_Y3.coord_z = 1;
defparam syncload_ctrl_X59_Y3.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X59_Y4(
	.Din(),
	.Dout(SyncLoad_X59_Y4_VCC));
defparam syncload_ctrl_X59_Y4.coord_x = 17;
defparam syncload_ctrl_X59_Y4.coord_y = 11;
defparam syncload_ctrl_X59_Y4.coord_z = 1;
defparam syncload_ctrl_X59_Y4.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X59_Y5(
	.Din(),
	.Dout(SyncLoad_X59_Y5_VCC));
defparam syncload_ctrl_X59_Y5.coord_x = 14;
defparam syncload_ctrl_X59_Y5.coord_y = 8;
defparam syncload_ctrl_X59_Y5.coord_z = 1;
defparam syncload_ctrl_X59_Y5.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X59_Y7(
	.Din(),
	.Dout(SyncLoad_X59_Y7_VCC));
defparam syncload_ctrl_X59_Y7.coord_x = 18;
defparam syncload_ctrl_X59_Y7.coord_y = 5;
defparam syncload_ctrl_X59_Y7.coord_z = 1;
defparam syncload_ctrl_X59_Y7.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X59_Y8(
	.Din(),
	.Dout(SyncLoad_X59_Y8_VCC));
defparam syncload_ctrl_X59_Y8.coord_x = 14;
defparam syncload_ctrl_X59_Y8.coord_y = 6;
defparam syncload_ctrl_X59_Y8.coord_z = 1;
defparam syncload_ctrl_X59_Y8.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X59_Y9(
	.Din(),
	.Dout(SyncLoad_X59_Y9_VCC));
defparam syncload_ctrl_X59_Y9.coord_x = 18;
defparam syncload_ctrl_X59_Y9.coord_y = 10;
defparam syncload_ctrl_X59_Y9.coord_z = 1;
defparam syncload_ctrl_X59_Y9.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X60_Y1(
	.Din(),
	.Dout(SyncLoad_X60_Y1_VCC));
defparam syncload_ctrl_X60_Y1.coord_x = 17;
defparam syncload_ctrl_X60_Y1.coord_y = 1;
defparam syncload_ctrl_X60_Y1.coord_z = 1;
defparam syncload_ctrl_X60_Y1.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X60_Y10(
	.Din(),
	.Dout(SyncLoad_X60_Y10_VCC));
defparam syncload_ctrl_X60_Y10.coord_x = 20;
defparam syncload_ctrl_X60_Y10.coord_y = 11;
defparam syncload_ctrl_X60_Y10.coord_z = 1;
defparam syncload_ctrl_X60_Y10.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X60_Y11(
	.Din(),
	.Dout(SyncLoad_X60_Y11_VCC));
defparam syncload_ctrl_X60_Y11.coord_x = 19;
defparam syncload_ctrl_X60_Y11.coord_y = 4;
defparam syncload_ctrl_X60_Y11.coord_z = 1;
defparam syncload_ctrl_X60_Y11.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X60_Y12(
	.Din(),
	.Dout(SyncLoad_X60_Y12_VCC));
defparam syncload_ctrl_X60_Y12.coord_x = 20;
defparam syncload_ctrl_X60_Y12.coord_y = 7;
defparam syncload_ctrl_X60_Y12.coord_z = 1;
defparam syncload_ctrl_X60_Y12.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X60_Y2(
	.Din(),
	.Dout(SyncLoad_X60_Y2_VCC));
defparam syncload_ctrl_X60_Y2.coord_x = 11;
defparam syncload_ctrl_X60_Y2.coord_y = 4;
defparam syncload_ctrl_X60_Y2.coord_z = 1;
defparam syncload_ctrl_X60_Y2.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X60_Y3(
	.Din(),
	.Dout(SyncLoad_X60_Y3_VCC));
defparam syncload_ctrl_X60_Y3.coord_x = 15;
defparam syncload_ctrl_X60_Y3.coord_y = 7;
defparam syncload_ctrl_X60_Y3.coord_z = 1;
defparam syncload_ctrl_X60_Y3.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X60_Y4(
	.Din(),
	.Dout(SyncLoad_X60_Y4_VCC));
defparam syncload_ctrl_X60_Y4.coord_x = 15;
defparam syncload_ctrl_X60_Y4.coord_y = 8;
defparam syncload_ctrl_X60_Y4.coord_z = 1;
defparam syncload_ctrl_X60_Y4.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X60_Y5(
	.Din(),
	.Dout(SyncLoad_X60_Y5_VCC));
defparam syncload_ctrl_X60_Y5.coord_x = 15;
defparam syncload_ctrl_X60_Y5.coord_y = 10;
defparam syncload_ctrl_X60_Y5.coord_z = 1;
defparam syncload_ctrl_X60_Y5.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X60_Y6(
	.Din(),
	.Dout(SyncLoad_X60_Y6_VCC));
defparam syncload_ctrl_X60_Y6.coord_x = 18;
defparam syncload_ctrl_X60_Y6.coord_y = 7;
defparam syncload_ctrl_X60_Y6.coord_z = 1;
defparam syncload_ctrl_X60_Y6.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X60_Y7(
	.Din(),
	.Dout(SyncLoad_X60_Y7_VCC));
defparam syncload_ctrl_X60_Y7.coord_x = 18;
defparam syncload_ctrl_X60_Y7.coord_y = 4;
defparam syncload_ctrl_X60_Y7.coord_z = 1;
defparam syncload_ctrl_X60_Y7.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X60_Y8(
	.Din(),
	.Dout(SyncLoad_X60_Y8_VCC));
defparam syncload_ctrl_X60_Y8.coord_x = 16;
defparam syncload_ctrl_X60_Y8.coord_y = 7;
defparam syncload_ctrl_X60_Y8.coord_z = 1;
defparam syncload_ctrl_X60_Y8.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X60_Y9(
	.Din(),
	.Dout(SyncLoad_X60_Y9_VCC));
defparam syncload_ctrl_X60_Y9.coord_x = 20;
defparam syncload_ctrl_X60_Y9.coord_y = 4;
defparam syncload_ctrl_X60_Y9.coord_z = 1;
defparam syncload_ctrl_X60_Y9.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X61_Y1(
	.Din(),
	.Dout(SyncLoad_X61_Y1_VCC));
defparam syncload_ctrl_X61_Y1.coord_x = 18;
defparam syncload_ctrl_X61_Y1.coord_y = 1;
defparam syncload_ctrl_X61_Y1.coord_z = 1;
defparam syncload_ctrl_X61_Y1.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X61_Y10(
	.Din(),
	.Dout(SyncLoad_X61_Y10_VCC));
defparam syncload_ctrl_X61_Y10.coord_x = 19;
defparam syncload_ctrl_X61_Y10.coord_y = 9;
defparam syncload_ctrl_X61_Y10.coord_z = 1;
defparam syncload_ctrl_X61_Y10.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X61_Y11(
	.Din(),
	.Dout(SyncLoad_X61_Y11_VCC));
defparam syncload_ctrl_X61_Y11.coord_x = 19;
defparam syncload_ctrl_X61_Y11.coord_y = 8;
defparam syncload_ctrl_X61_Y11.coord_z = 1;
defparam syncload_ctrl_X61_Y11.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X61_Y2(
	.Din(),
	.Dout(SyncLoad_X61_Y2_VCC));
defparam syncload_ctrl_X61_Y2.coord_x = 15;
defparam syncload_ctrl_X61_Y2.coord_y = 5;
defparam syncload_ctrl_X61_Y2.coord_z = 1;
defparam syncload_ctrl_X61_Y2.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X61_Y3(
	.Din(),
	.Dout(SyncLoad_X61_Y3_VCC));
defparam syncload_ctrl_X61_Y3.coord_x = 15;
defparam syncload_ctrl_X61_Y3.coord_y = 1;
defparam syncload_ctrl_X61_Y3.coord_z = 1;
defparam syncload_ctrl_X61_Y3.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X61_Y4(
	.Din(),
	.Dout(SyncLoad_X61_Y4_VCC));
defparam syncload_ctrl_X61_Y4.coord_x = 17;
defparam syncload_ctrl_X61_Y4.coord_y = 8;
defparam syncload_ctrl_X61_Y4.coord_z = 1;
defparam syncload_ctrl_X61_Y4.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X61_Y5(
	.Din(),
	.Dout(SyncLoad_X61_Y5_VCC));
defparam syncload_ctrl_X61_Y5.coord_x = 14;
defparam syncload_ctrl_X61_Y5.coord_y = 1;
defparam syncload_ctrl_X61_Y5.coord_z = 1;
defparam syncload_ctrl_X61_Y5.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X61_Y6(
	.Din(),
	.Dout(SyncLoad_X61_Y6_VCC));
defparam syncload_ctrl_X61_Y6.coord_x = 15;
defparam syncload_ctrl_X61_Y6.coord_y = 9;
defparam syncload_ctrl_X61_Y6.coord_z = 1;
defparam syncload_ctrl_X61_Y6.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X61_Y7(
	.Din(),
	.Dout(SyncLoad_X61_Y7_VCC));
defparam syncload_ctrl_X61_Y7.coord_x = 17;
defparam syncload_ctrl_X61_Y7.coord_y = 3;
defparam syncload_ctrl_X61_Y7.coord_z = 1;
defparam syncload_ctrl_X61_Y7.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X61_Y8(
	.Din(),
	.Dout(SyncLoad_X61_Y8_VCC));
defparam syncload_ctrl_X61_Y8.coord_x = 19;
defparam syncload_ctrl_X61_Y8.coord_y = 2;
defparam syncload_ctrl_X61_Y8.coord_z = 1;
defparam syncload_ctrl_X61_Y8.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X61_Y9(
	.Din(),
	.Dout(SyncLoad_X61_Y9_VCC));
defparam syncload_ctrl_X61_Y9.coord_x = 19;
defparam syncload_ctrl_X61_Y9.coord_y = 7;
defparam syncload_ctrl_X61_Y9.coord_z = 1;
defparam syncload_ctrl_X61_Y9.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X62_Y1(
	.Din(),
	.Dout(SyncLoad_X62_Y1_VCC));
defparam syncload_ctrl_X62_Y1.coord_x = 12;
defparam syncload_ctrl_X62_Y1.coord_y = 1;
defparam syncload_ctrl_X62_Y1.coord_z = 1;
defparam syncload_ctrl_X62_Y1.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X62_Y10(
	.Din(),
	.Dout(SyncLoad_X62_Y10_VCC));
defparam syncload_ctrl_X62_Y10.coord_x = 20;
defparam syncload_ctrl_X62_Y10.coord_y = 12;
defparam syncload_ctrl_X62_Y10.coord_z = 1;
defparam syncload_ctrl_X62_Y10.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X62_Y11(
	.Din(),
	.Dout(SyncLoad_X62_Y11_VCC));
defparam syncload_ctrl_X62_Y11.coord_x = 20;
defparam syncload_ctrl_X62_Y11.coord_y = 9;
defparam syncload_ctrl_X62_Y11.coord_z = 1;
defparam syncload_ctrl_X62_Y11.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X62_Y2(
	.Din(),
	.Dout(SyncLoad_X62_Y2_VCC));
defparam syncload_ctrl_X62_Y2.coord_x = 17;
defparam syncload_ctrl_X62_Y2.coord_y = 6;
defparam syncload_ctrl_X62_Y2.coord_z = 1;
defparam syncload_ctrl_X62_Y2.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X62_Y3(
	.Din(),
	.Dout(SyncLoad_X62_Y3_VCC));
defparam syncload_ctrl_X62_Y3.coord_x = 16;
defparam syncload_ctrl_X62_Y3.coord_y = 6;
defparam syncload_ctrl_X62_Y3.coord_z = 1;
defparam syncload_ctrl_X62_Y3.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X62_Y4(
	.Din(),
	.Dout(SyncLoad_X62_Y4_VCC));
defparam syncload_ctrl_X62_Y4.coord_x = 14;
defparam syncload_ctrl_X62_Y4.coord_y = 3;
defparam syncload_ctrl_X62_Y4.coord_z = 1;
defparam syncload_ctrl_X62_Y4.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X62_Y5(
	.Din(),
	.Dout(SyncLoad_X62_Y5_VCC));
defparam syncload_ctrl_X62_Y5.coord_x = 17;
defparam syncload_ctrl_X62_Y5.coord_y = 10;
defparam syncload_ctrl_X62_Y5.coord_z = 1;
defparam syncload_ctrl_X62_Y5.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X62_Y6(
	.Din(),
	.Dout(SyncLoad_X62_Y6_VCC));
defparam syncload_ctrl_X62_Y6.coord_x = 17;
defparam syncload_ctrl_X62_Y6.coord_y = 12;
defparam syncload_ctrl_X62_Y6.coord_z = 1;
defparam syncload_ctrl_X62_Y6.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X62_Y7(
	.Din(),
	.Dout(SyncLoad_X62_Y7_VCC));
defparam syncload_ctrl_X62_Y7.coord_x = 15;
defparam syncload_ctrl_X62_Y7.coord_y = 6;
defparam syncload_ctrl_X62_Y7.coord_z = 1;
defparam syncload_ctrl_X62_Y7.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X62_Y8(
	.Din(),
	.Dout(SyncLoad_X62_Y8_VCC));
defparam syncload_ctrl_X62_Y8.coord_x = 18;
defparam syncload_ctrl_X62_Y8.coord_y = 2;
defparam syncload_ctrl_X62_Y8.coord_z = 1;
defparam syncload_ctrl_X62_Y8.SyncCtrlMux = 2'b01;

alta_syncctrl syncload_ctrl_X62_Y9(
	.Din(),
	.Dout(SyncLoad_X62_Y9_VCC));
defparam syncload_ctrl_X62_Y9.coord_x = 19;
defparam syncload_ctrl_X62_Y9.coord_y = 11;
defparam syncload_ctrl_X62_Y9.coord_z = 1;
defparam syncload_ctrl_X62_Y9.SyncCtrlMux = 2'b01;

alta_syncctrl syncreset_ctrl_X43_Y2(
	.Din(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout ),
	.Dout(\macro_inst|serial_lim_input_inst|shift_div_counter[2]~20_combout__SyncReset_X43_Y2_SIG ));
defparam syncreset_ctrl_X43_Y2.coord_x = 7;
defparam syncreset_ctrl_X43_Y2.coord_y = 2;
defparam syncreset_ctrl_X43_Y2.coord_z = 0;
defparam syncreset_ctrl_X43_Y2.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X46_Y2(
	.Din(),
	.Dout(SyncReset_X46_Y2_GND));
defparam syncreset_ctrl_X46_Y2.coord_x = 4;
defparam syncreset_ctrl_X46_Y2.coord_y = 3;
defparam syncreset_ctrl_X46_Y2.coord_z = 0;
defparam syncreset_ctrl_X46_Y2.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X46_Y3(
	.Din(),
	.Dout(SyncReset_X46_Y3_GND));
defparam syncreset_ctrl_X46_Y3.coord_x = 5;
defparam syncreset_ctrl_X46_Y3.coord_y = 4;
defparam syncreset_ctrl_X46_Y3.coord_z = 0;
defparam syncreset_ctrl_X46_Y3.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X47_Y3(
	.Din(),
	.Dout(SyncReset_X47_Y3_GND));
defparam syncreset_ctrl_X47_Y3.coord_x = 4;
defparam syncreset_ctrl_X47_Y3.coord_y = 4;
defparam syncreset_ctrl_X47_Y3.coord_z = 0;
defparam syncreset_ctrl_X47_Y3.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X49_Y2(
	.Din(),
	.Dout(SyncReset_X49_Y2_GND));
defparam syncreset_ctrl_X49_Y2.coord_x = 9;
defparam syncreset_ctrl_X49_Y2.coord_y = 3;
defparam syncreset_ctrl_X49_Y2.coord_z = 0;
defparam syncreset_ctrl_X49_Y2.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X49_Y3(
	.Din(),
	.Dout(SyncReset_X49_Y3_GND));
defparam syncreset_ctrl_X49_Y3.coord_x = 6;
defparam syncreset_ctrl_X49_Y3.coord_y = 4;
defparam syncreset_ctrl_X49_Y3.coord_z = 0;
defparam syncreset_ctrl_X49_Y3.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X50_Y1(
	.Din(),
	.Dout(SyncReset_X50_Y1_GND));
defparam syncreset_ctrl_X50_Y1.coord_x = 7;
defparam syncreset_ctrl_X50_Y1.coord_y = 1;
defparam syncreset_ctrl_X50_Y1.coord_z = 0;
defparam syncreset_ctrl_X50_Y1.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X50_Y2(
	.Din(\macro_inst|controller|serial|bit_counter[7]~17_combout ),
	.Dout(\macro_inst|controller|serial|bit_counter[7]~17_combout__SyncReset_X50_Y2_SIG ));
defparam syncreset_ctrl_X50_Y2.coord_x = 9;
defparam syncreset_ctrl_X50_Y2.coord_y = 2;
defparam syncreset_ctrl_X50_Y2.coord_z = 0;
defparam syncreset_ctrl_X50_Y2.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X50_Y3(
	.Din(),
	.Dout(SyncReset_X50_Y3_GND));
defparam syncreset_ctrl_X50_Y3.coord_x = 8;
defparam syncreset_ctrl_X50_Y3.coord_y = 4;
defparam syncreset_ctrl_X50_Y3.coord_z = 0;
defparam syncreset_ctrl_X50_Y3.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X51_Y2(
	.Din(\macro_inst|controller|serial|state.IDLE~q ),
	.Dout(\macro_inst|controller|serial|state.IDLE~q__SyncReset_X51_Y2_INV ));
defparam syncreset_ctrl_X51_Y2.coord_x = 8;
defparam syncreset_ctrl_X51_Y2.coord_y = 2;
defparam syncreset_ctrl_X51_Y2.coord_z = 0;
defparam syncreset_ctrl_X51_Y2.SyncCtrlMux = 2'b11;

alta_syncctrl syncreset_ctrl_X51_Y3(
	.Din(),
	.Dout(SyncReset_X51_Y3_GND));
defparam syncreset_ctrl_X51_Y3.coord_x = 9;
defparam syncreset_ctrl_X51_Y3.coord_y = 4;
defparam syncreset_ctrl_X51_Y3.coord_z = 0;
defparam syncreset_ctrl_X51_Y3.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X51_Y4(
	.Din(),
	.Dout(SyncReset_X51_Y4_GND));
defparam syncreset_ctrl_X51_Y4.coord_x = 15;
defparam syncreset_ctrl_X51_Y4.coord_y = 2;
defparam syncreset_ctrl_X51_Y4.coord_z = 0;
defparam syncreset_ctrl_X51_Y4.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X52_Y2(
	.Din(),
	.Dout(SyncReset_X52_Y2_GND));
defparam syncreset_ctrl_X52_Y2.coord_x = 16;
defparam syncreset_ctrl_X52_Y2.coord_y = 5;
defparam syncreset_ctrl_X52_Y2.coord_z = 0;
defparam syncreset_ctrl_X52_Y2.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X52_Y3(
	.Din(),
	.Dout(SyncReset_X52_Y3_GND));
defparam syncreset_ctrl_X52_Y3.coord_x = 8;
defparam syncreset_ctrl_X52_Y3.coord_y = 3;
defparam syncreset_ctrl_X52_Y3.coord_z = 0;
defparam syncreset_ctrl_X52_Y3.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X52_Y4(
	.Din(),
	.Dout(SyncReset_X52_Y4_GND));
defparam syncreset_ctrl_X52_Y4.coord_x = 16;
defparam syncreset_ctrl_X52_Y4.coord_y = 2;
defparam syncreset_ctrl_X52_Y4.coord_z = 0;
defparam syncreset_ctrl_X52_Y4.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X53_Y4(
	.Din(),
	.Dout(SyncReset_X53_Y4_GND));
defparam syncreset_ctrl_X53_Y4.coord_x = 15;
defparam syncreset_ctrl_X53_Y4.coord_y = 4;
defparam syncreset_ctrl_X53_Y4.coord_z = 0;
defparam syncreset_ctrl_X53_Y4.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X54_Y1(
	.Din(),
	.Dout(SyncReset_X54_Y1_GND));
defparam syncreset_ctrl_X54_Y1.coord_x = 20;
defparam syncreset_ctrl_X54_Y1.coord_y = 2;
defparam syncreset_ctrl_X54_Y1.coord_z = 0;
defparam syncreset_ctrl_X54_Y1.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X54_Y2(
	.Din(),
	.Dout(SyncReset_X54_Y2_GND));
defparam syncreset_ctrl_X54_Y2.coord_x = 14;
defparam syncreset_ctrl_X54_Y2.coord_y = 5;
defparam syncreset_ctrl_X54_Y2.coord_z = 0;
defparam syncreset_ctrl_X54_Y2.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X54_Y3(
	.Din(),
	.Dout(SyncReset_X54_Y3_GND));
defparam syncreset_ctrl_X54_Y3.coord_x = 14;
defparam syncreset_ctrl_X54_Y3.coord_y = 12;
defparam syncreset_ctrl_X54_Y3.coord_z = 0;
defparam syncreset_ctrl_X54_Y3.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X54_Y4(
	.Din(),
	.Dout(SyncReset_X54_Y4_GND));
defparam syncreset_ctrl_X54_Y4.coord_x = 11;
defparam syncreset_ctrl_X54_Y4.coord_y = 2;
defparam syncreset_ctrl_X54_Y4.coord_z = 0;
defparam syncreset_ctrl_X54_Y4.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X56_Y1(
	.Din(),
	.Dout(SyncReset_X56_Y1_GND));
defparam syncreset_ctrl_X56_Y1.coord_x = 10;
defparam syncreset_ctrl_X56_Y1.coord_y = 2;
defparam syncreset_ctrl_X56_Y1.coord_z = 0;
defparam syncreset_ctrl_X56_Y1.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X56_Y10(
	.Din(),
	.Dout(SyncReset_X56_Y10_GND));
defparam syncreset_ctrl_X56_Y10.coord_x = 11;
defparam syncreset_ctrl_X56_Y10.coord_y = 3;
defparam syncreset_ctrl_X56_Y10.coord_z = 0;
defparam syncreset_ctrl_X56_Y10.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X56_Y2(
	.Din(),
	.Dout(SyncReset_X56_Y2_GND));
defparam syncreset_ctrl_X56_Y2.coord_x = 16;
defparam syncreset_ctrl_X56_Y2.coord_y = 11;
defparam syncreset_ctrl_X56_Y2.coord_z = 0;
defparam syncreset_ctrl_X56_Y2.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X56_Y3(
	.Din(\rv32.mem_ahb_haddr[3] ),
	.Dout(\rv32.mem_ahb_haddr[3]__SyncReset_X56_Y3_SIG ));
defparam syncreset_ctrl_X56_Y3.coord_x = 12;
defparam syncreset_ctrl_X56_Y3.coord_y = 4;
defparam syncreset_ctrl_X56_Y3.coord_z = 0;
defparam syncreset_ctrl_X56_Y3.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X56_Y4(
	.Din(),
	.Dout(SyncReset_X56_Y4_GND));
defparam syncreset_ctrl_X56_Y4.coord_x = 17;
defparam syncreset_ctrl_X56_Y4.coord_y = 4;
defparam syncreset_ctrl_X56_Y4.coord_z = 0;
defparam syncreset_ctrl_X56_Y4.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X56_Y5(
	.Din(\rv32.mem_ahb_haddr[3] ),
	.Dout(\rv32.mem_ahb_haddr[3]__SyncReset_X56_Y5_SIG ));
defparam syncreset_ctrl_X56_Y5.coord_x = 10;
defparam syncreset_ctrl_X56_Y5.coord_y = 4;
defparam syncreset_ctrl_X56_Y5.coord_z = 0;
defparam syncreset_ctrl_X56_Y5.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X56_Y6(
	.Din(),
	.Dout(SyncReset_X56_Y6_GND));
defparam syncreset_ctrl_X56_Y6.coord_x = 17;
defparam syncreset_ctrl_X56_Y6.coord_y = 2;
defparam syncreset_ctrl_X56_Y6.coord_z = 0;
defparam syncreset_ctrl_X56_Y6.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X56_Y7(
	.Din(),
	.Dout(SyncReset_X56_Y7_GND));
defparam syncreset_ctrl_X56_Y7.coord_x = 14;
defparam syncreset_ctrl_X56_Y7.coord_y = 2;
defparam syncreset_ctrl_X56_Y7.coord_z = 0;
defparam syncreset_ctrl_X56_Y7.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X56_Y8(
	.Din(),
	.Dout(SyncReset_X56_Y8_GND));
defparam syncreset_ctrl_X56_Y8.coord_x = 19;
defparam syncreset_ctrl_X56_Y8.coord_y = 1;
defparam syncreset_ctrl_X56_Y8.coord_z = 0;
defparam syncreset_ctrl_X56_Y8.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X56_Y9(
	.Din(),
	.Dout(SyncReset_X56_Y9_GND));
defparam syncreset_ctrl_X56_Y9.coord_x = 17;
defparam syncreset_ctrl_X56_Y9.coord_y = 9;
defparam syncreset_ctrl_X56_Y9.coord_z = 0;
defparam syncreset_ctrl_X56_Y9.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X57_Y1(
	.Din(),
	.Dout(SyncReset_X57_Y1_GND));
defparam syncreset_ctrl_X57_Y1.coord_x = 12;
defparam syncreset_ctrl_X57_Y1.coord_y = 2;
defparam syncreset_ctrl_X57_Y1.coord_z = 0;
defparam syncreset_ctrl_X57_Y1.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X57_Y10(
	.Din(),
	.Dout(SyncReset_X57_Y10_GND));
defparam syncreset_ctrl_X57_Y10.coord_x = 12;
defparam syncreset_ctrl_X57_Y10.coord_y = 3;
defparam syncreset_ctrl_X57_Y10.coord_z = 0;
defparam syncreset_ctrl_X57_Y10.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X57_Y11(
	.Din(),
	.Dout(SyncReset_X57_Y11_GND));
defparam syncreset_ctrl_X57_Y11.coord_x = 20;
defparam syncreset_ctrl_X57_Y11.coord_y = 10;
defparam syncreset_ctrl_X57_Y11.coord_z = 0;
defparam syncreset_ctrl_X57_Y11.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X57_Y12(
	.Din(),
	.Dout(SyncReset_X57_Y12_GND));
defparam syncreset_ctrl_X57_Y12.coord_x = 18;
defparam syncreset_ctrl_X57_Y12.coord_y = 8;
defparam syncreset_ctrl_X57_Y12.coord_z = 0;
defparam syncreset_ctrl_X57_Y12.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X57_Y2(
	.Din(),
	.Dout(SyncReset_X57_Y2_GND));
defparam syncreset_ctrl_X57_Y2.coord_x = 18;
defparam syncreset_ctrl_X57_Y2.coord_y = 12;
defparam syncreset_ctrl_X57_Y2.coord_z = 0;
defparam syncreset_ctrl_X57_Y2.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X57_Y3(
	.Din(),
	.Dout(SyncReset_X57_Y3_GND));
defparam syncreset_ctrl_X57_Y3.coord_x = 14;
defparam syncreset_ctrl_X57_Y3.coord_y = 11;
defparam syncreset_ctrl_X57_Y3.coord_z = 0;
defparam syncreset_ctrl_X57_Y3.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X57_Y4(
	.Din(),
	.Dout(SyncReset_X57_Y4_GND));
defparam syncreset_ctrl_X57_Y4.coord_x = 16;
defparam syncreset_ctrl_X57_Y4.coord_y = 4;
defparam syncreset_ctrl_X57_Y4.coord_z = 0;
defparam syncreset_ctrl_X57_Y4.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X57_Y5(
	.Din(\rv32.mem_ahb_haddr[3] ),
	.Dout(\rv32.mem_ahb_haddr[3]__SyncReset_X57_Y5_SIG ));
defparam syncreset_ctrl_X57_Y5.coord_x = 14;
defparam syncreset_ctrl_X57_Y5.coord_y = 7;
defparam syncreset_ctrl_X57_Y5.coord_z = 0;
defparam syncreset_ctrl_X57_Y5.SyncCtrlMux = 2'b10;

alta_syncctrl syncreset_ctrl_X57_Y6(
	.Din(),
	.Dout(SyncReset_X57_Y6_GND));
defparam syncreset_ctrl_X57_Y6.coord_x = 14;
defparam syncreset_ctrl_X57_Y6.coord_y = 10;
defparam syncreset_ctrl_X57_Y6.coord_z = 0;
defparam syncreset_ctrl_X57_Y6.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X57_Y8(
	.Din(),
	.Dout(SyncReset_X57_Y8_GND));
defparam syncreset_ctrl_X57_Y8.coord_x = 18;
defparam syncreset_ctrl_X57_Y8.coord_y = 3;
defparam syncreset_ctrl_X57_Y8.coord_z = 0;
defparam syncreset_ctrl_X57_Y8.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X57_Y9(
	.Din(),
	.Dout(SyncReset_X57_Y9_GND));
defparam syncreset_ctrl_X57_Y9.coord_x = 16;
defparam syncreset_ctrl_X57_Y9.coord_y = 9;
defparam syncreset_ctrl_X57_Y9.coord_z = 0;
defparam syncreset_ctrl_X57_Y9.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X58_Y1(
	.Din(),
	.Dout(SyncReset_X58_Y1_GND));
defparam syncreset_ctrl_X58_Y1.coord_x = 10;
defparam syncreset_ctrl_X58_Y1.coord_y = 1;
defparam syncreset_ctrl_X58_Y1.coord_z = 0;
defparam syncreset_ctrl_X58_Y1.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X58_Y10(
	.Din(),
	.Dout(SyncReset_X58_Y10_GND));
defparam syncreset_ctrl_X58_Y10.coord_x = 17;
defparam syncreset_ctrl_X58_Y10.coord_y = 7;
defparam syncreset_ctrl_X58_Y10.coord_z = 0;
defparam syncreset_ctrl_X58_Y10.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X58_Y11(
	.Din(),
	.Dout(SyncReset_X58_Y11_GND));
defparam syncreset_ctrl_X58_Y11.coord_x = 19;
defparam syncreset_ctrl_X58_Y11.coord_y = 12;
defparam syncreset_ctrl_X58_Y11.coord_z = 0;
defparam syncreset_ctrl_X58_Y11.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X58_Y12(
	.Din(),
	.Dout(SyncReset_X58_Y12_GND));
defparam syncreset_ctrl_X58_Y12.coord_x = 20;
defparam syncreset_ctrl_X58_Y12.coord_y = 3;
defparam syncreset_ctrl_X58_Y12.coord_z = 0;
defparam syncreset_ctrl_X58_Y12.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X58_Y2(
	.Din(),
	.Dout(SyncReset_X58_Y2_GND));
defparam syncreset_ctrl_X58_Y2.coord_x = 16;
defparam syncreset_ctrl_X58_Y2.coord_y = 10;
defparam syncreset_ctrl_X58_Y2.coord_z = 0;
defparam syncreset_ctrl_X58_Y2.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X58_Y3(
	.Din(),
	.Dout(SyncReset_X58_Y3_GND));
defparam syncreset_ctrl_X58_Y3.coord_x = 15;
defparam syncreset_ctrl_X58_Y3.coord_y = 11;
defparam syncreset_ctrl_X58_Y3.coord_z = 0;
defparam syncreset_ctrl_X58_Y3.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X58_Y4(
	.Din(),
	.Dout(SyncReset_X58_Y4_GND));
defparam syncreset_ctrl_X58_Y4.coord_x = 16;
defparam syncreset_ctrl_X58_Y4.coord_y = 8;
defparam syncreset_ctrl_X58_Y4.coord_z = 0;
defparam syncreset_ctrl_X58_Y4.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X58_Y5(
	.Din(),
	.Dout(SyncReset_X58_Y5_GND));
defparam syncreset_ctrl_X58_Y5.coord_x = 16;
defparam syncreset_ctrl_X58_Y5.coord_y = 12;
defparam syncreset_ctrl_X58_Y5.coord_z = 0;
defparam syncreset_ctrl_X58_Y5.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X58_Y6(
	.Din(),
	.Dout(SyncReset_X58_Y6_GND));
defparam syncreset_ctrl_X58_Y6.coord_x = 14;
defparam syncreset_ctrl_X58_Y6.coord_y = 9;
defparam syncreset_ctrl_X58_Y6.coord_z = 0;
defparam syncreset_ctrl_X58_Y6.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X58_Y7(
	.Din(),
	.Dout(SyncReset_X58_Y7_GND));
defparam syncreset_ctrl_X58_Y7.coord_x = 14;
defparam syncreset_ctrl_X58_Y7.coord_y = 4;
defparam syncreset_ctrl_X58_Y7.coord_z = 0;
defparam syncreset_ctrl_X58_Y7.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X58_Y8(
	.Din(),
	.Dout(SyncReset_X58_Y8_GND));
defparam syncreset_ctrl_X58_Y8.coord_x = 17;
defparam syncreset_ctrl_X58_Y8.coord_y = 5;
defparam syncreset_ctrl_X58_Y8.coord_z = 0;
defparam syncreset_ctrl_X58_Y8.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X58_Y9(
	.Din(),
	.Dout(SyncReset_X58_Y9_GND));
defparam syncreset_ctrl_X58_Y9.coord_x = 18;
defparam syncreset_ctrl_X58_Y9.coord_y = 9;
defparam syncreset_ctrl_X58_Y9.coord_z = 0;
defparam syncreset_ctrl_X58_Y9.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X59_Y1(
	.Din(),
	.Dout(SyncReset_X59_Y1_GND));
defparam syncreset_ctrl_X59_Y1.coord_x = 16;
defparam syncreset_ctrl_X59_Y1.coord_y = 3;
defparam syncreset_ctrl_X59_Y1.coord_z = 0;
defparam syncreset_ctrl_X59_Y1.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X59_Y10(
	.Din(),
	.Dout(SyncReset_X59_Y10_GND));
defparam syncreset_ctrl_X59_Y10.coord_x = 18;
defparam syncreset_ctrl_X59_Y10.coord_y = 6;
defparam syncreset_ctrl_X59_Y10.coord_z = 0;
defparam syncreset_ctrl_X59_Y10.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X59_Y11(
	.Din(),
	.Dout(SyncReset_X59_Y11_GND));
defparam syncreset_ctrl_X59_Y11.coord_x = 19;
defparam syncreset_ctrl_X59_Y11.coord_y = 3;
defparam syncreset_ctrl_X59_Y11.coord_z = 0;
defparam syncreset_ctrl_X59_Y11.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X59_Y12(
	.Din(),
	.Dout(SyncReset_X59_Y12_GND));
defparam syncreset_ctrl_X59_Y12.coord_x = 20;
defparam syncreset_ctrl_X59_Y12.coord_y = 5;
defparam syncreset_ctrl_X59_Y12.coord_z = 0;
defparam syncreset_ctrl_X59_Y12.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X59_Y2(
	.Din(),
	.Dout(SyncReset_X59_Y2_GND));
defparam syncreset_ctrl_X59_Y2.coord_x = 10;
defparam syncreset_ctrl_X59_Y2.coord_y = 3;
defparam syncreset_ctrl_X59_Y2.coord_z = 0;
defparam syncreset_ctrl_X59_Y2.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X59_Y3(
	.Din(),
	.Dout(SyncReset_X59_Y3_GND));
defparam syncreset_ctrl_X59_Y3.coord_x = 15;
defparam syncreset_ctrl_X59_Y3.coord_y = 12;
defparam syncreset_ctrl_X59_Y3.coord_z = 0;
defparam syncreset_ctrl_X59_Y3.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X59_Y4(
	.Din(),
	.Dout(SyncReset_X59_Y4_GND));
defparam syncreset_ctrl_X59_Y4.coord_x = 17;
defparam syncreset_ctrl_X59_Y4.coord_y = 11;
defparam syncreset_ctrl_X59_Y4.coord_z = 0;
defparam syncreset_ctrl_X59_Y4.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X59_Y5(
	.Din(),
	.Dout(SyncReset_X59_Y5_GND));
defparam syncreset_ctrl_X59_Y5.coord_x = 14;
defparam syncreset_ctrl_X59_Y5.coord_y = 8;
defparam syncreset_ctrl_X59_Y5.coord_z = 0;
defparam syncreset_ctrl_X59_Y5.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X59_Y7(
	.Din(),
	.Dout(SyncReset_X59_Y7_GND));
defparam syncreset_ctrl_X59_Y7.coord_x = 18;
defparam syncreset_ctrl_X59_Y7.coord_y = 5;
defparam syncreset_ctrl_X59_Y7.coord_z = 0;
defparam syncreset_ctrl_X59_Y7.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X59_Y8(
	.Din(),
	.Dout(SyncReset_X59_Y8_GND));
defparam syncreset_ctrl_X59_Y8.coord_x = 14;
defparam syncreset_ctrl_X59_Y8.coord_y = 6;
defparam syncreset_ctrl_X59_Y8.coord_z = 0;
defparam syncreset_ctrl_X59_Y8.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X59_Y9(
	.Din(),
	.Dout(SyncReset_X59_Y9_GND));
defparam syncreset_ctrl_X59_Y9.coord_x = 18;
defparam syncreset_ctrl_X59_Y9.coord_y = 10;
defparam syncreset_ctrl_X59_Y9.coord_z = 0;
defparam syncreset_ctrl_X59_Y9.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X60_Y1(
	.Din(),
	.Dout(SyncReset_X60_Y1_GND));
defparam syncreset_ctrl_X60_Y1.coord_x = 17;
defparam syncreset_ctrl_X60_Y1.coord_y = 1;
defparam syncreset_ctrl_X60_Y1.coord_z = 0;
defparam syncreset_ctrl_X60_Y1.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X60_Y10(
	.Din(),
	.Dout(SyncReset_X60_Y10_GND));
defparam syncreset_ctrl_X60_Y10.coord_x = 20;
defparam syncreset_ctrl_X60_Y10.coord_y = 11;
defparam syncreset_ctrl_X60_Y10.coord_z = 0;
defparam syncreset_ctrl_X60_Y10.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X60_Y11(
	.Din(),
	.Dout(SyncReset_X60_Y11_GND));
defparam syncreset_ctrl_X60_Y11.coord_x = 19;
defparam syncreset_ctrl_X60_Y11.coord_y = 4;
defparam syncreset_ctrl_X60_Y11.coord_z = 0;
defparam syncreset_ctrl_X60_Y11.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X60_Y12(
	.Din(),
	.Dout(SyncReset_X60_Y12_GND));
defparam syncreset_ctrl_X60_Y12.coord_x = 20;
defparam syncreset_ctrl_X60_Y12.coord_y = 7;
defparam syncreset_ctrl_X60_Y12.coord_z = 0;
defparam syncreset_ctrl_X60_Y12.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X60_Y2(
	.Din(),
	.Dout(SyncReset_X60_Y2_GND));
defparam syncreset_ctrl_X60_Y2.coord_x = 11;
defparam syncreset_ctrl_X60_Y2.coord_y = 4;
defparam syncreset_ctrl_X60_Y2.coord_z = 0;
defparam syncreset_ctrl_X60_Y2.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X60_Y3(
	.Din(),
	.Dout(SyncReset_X60_Y3_GND));
defparam syncreset_ctrl_X60_Y3.coord_x = 15;
defparam syncreset_ctrl_X60_Y3.coord_y = 7;
defparam syncreset_ctrl_X60_Y3.coord_z = 0;
defparam syncreset_ctrl_X60_Y3.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X60_Y4(
	.Din(),
	.Dout(SyncReset_X60_Y4_GND));
defparam syncreset_ctrl_X60_Y4.coord_x = 15;
defparam syncreset_ctrl_X60_Y4.coord_y = 8;
defparam syncreset_ctrl_X60_Y4.coord_z = 0;
defparam syncreset_ctrl_X60_Y4.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X60_Y5(
	.Din(),
	.Dout(SyncReset_X60_Y5_GND));
defparam syncreset_ctrl_X60_Y5.coord_x = 15;
defparam syncreset_ctrl_X60_Y5.coord_y = 10;
defparam syncreset_ctrl_X60_Y5.coord_z = 0;
defparam syncreset_ctrl_X60_Y5.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X60_Y6(
	.Din(),
	.Dout(SyncReset_X60_Y6_GND));
defparam syncreset_ctrl_X60_Y6.coord_x = 18;
defparam syncreset_ctrl_X60_Y6.coord_y = 7;
defparam syncreset_ctrl_X60_Y6.coord_z = 0;
defparam syncreset_ctrl_X60_Y6.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X60_Y7(
	.Din(),
	.Dout(SyncReset_X60_Y7_GND));
defparam syncreset_ctrl_X60_Y7.coord_x = 18;
defparam syncreset_ctrl_X60_Y7.coord_y = 4;
defparam syncreset_ctrl_X60_Y7.coord_z = 0;
defparam syncreset_ctrl_X60_Y7.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X60_Y8(
	.Din(),
	.Dout(SyncReset_X60_Y8_GND));
defparam syncreset_ctrl_X60_Y8.coord_x = 16;
defparam syncreset_ctrl_X60_Y8.coord_y = 7;
defparam syncreset_ctrl_X60_Y8.coord_z = 0;
defparam syncreset_ctrl_X60_Y8.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X60_Y9(
	.Din(),
	.Dout(SyncReset_X60_Y9_GND));
defparam syncreset_ctrl_X60_Y9.coord_x = 20;
defparam syncreset_ctrl_X60_Y9.coord_y = 4;
defparam syncreset_ctrl_X60_Y9.coord_z = 0;
defparam syncreset_ctrl_X60_Y9.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X61_Y1(
	.Din(),
	.Dout(SyncReset_X61_Y1_GND));
defparam syncreset_ctrl_X61_Y1.coord_x = 18;
defparam syncreset_ctrl_X61_Y1.coord_y = 1;
defparam syncreset_ctrl_X61_Y1.coord_z = 0;
defparam syncreset_ctrl_X61_Y1.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X61_Y10(
	.Din(),
	.Dout(SyncReset_X61_Y10_GND));
defparam syncreset_ctrl_X61_Y10.coord_x = 19;
defparam syncreset_ctrl_X61_Y10.coord_y = 9;
defparam syncreset_ctrl_X61_Y10.coord_z = 0;
defparam syncreset_ctrl_X61_Y10.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X61_Y11(
	.Din(),
	.Dout(SyncReset_X61_Y11_GND));
defparam syncreset_ctrl_X61_Y11.coord_x = 19;
defparam syncreset_ctrl_X61_Y11.coord_y = 8;
defparam syncreset_ctrl_X61_Y11.coord_z = 0;
defparam syncreset_ctrl_X61_Y11.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X61_Y2(
	.Din(),
	.Dout(SyncReset_X61_Y2_GND));
defparam syncreset_ctrl_X61_Y2.coord_x = 15;
defparam syncreset_ctrl_X61_Y2.coord_y = 5;
defparam syncreset_ctrl_X61_Y2.coord_z = 0;
defparam syncreset_ctrl_X61_Y2.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X61_Y3(
	.Din(),
	.Dout(SyncReset_X61_Y3_GND));
defparam syncreset_ctrl_X61_Y3.coord_x = 15;
defparam syncreset_ctrl_X61_Y3.coord_y = 1;
defparam syncreset_ctrl_X61_Y3.coord_z = 0;
defparam syncreset_ctrl_X61_Y3.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X61_Y4(
	.Din(),
	.Dout(SyncReset_X61_Y4_GND));
defparam syncreset_ctrl_X61_Y4.coord_x = 17;
defparam syncreset_ctrl_X61_Y4.coord_y = 8;
defparam syncreset_ctrl_X61_Y4.coord_z = 0;
defparam syncreset_ctrl_X61_Y4.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X61_Y5(
	.Din(),
	.Dout(SyncReset_X61_Y5_GND));
defparam syncreset_ctrl_X61_Y5.coord_x = 14;
defparam syncreset_ctrl_X61_Y5.coord_y = 1;
defparam syncreset_ctrl_X61_Y5.coord_z = 0;
defparam syncreset_ctrl_X61_Y5.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X61_Y6(
	.Din(),
	.Dout(SyncReset_X61_Y6_GND));
defparam syncreset_ctrl_X61_Y6.coord_x = 15;
defparam syncreset_ctrl_X61_Y6.coord_y = 9;
defparam syncreset_ctrl_X61_Y6.coord_z = 0;
defparam syncreset_ctrl_X61_Y6.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X61_Y7(
	.Din(),
	.Dout(SyncReset_X61_Y7_GND));
defparam syncreset_ctrl_X61_Y7.coord_x = 17;
defparam syncreset_ctrl_X61_Y7.coord_y = 3;
defparam syncreset_ctrl_X61_Y7.coord_z = 0;
defparam syncreset_ctrl_X61_Y7.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X61_Y8(
	.Din(),
	.Dout(SyncReset_X61_Y8_GND));
defparam syncreset_ctrl_X61_Y8.coord_x = 19;
defparam syncreset_ctrl_X61_Y8.coord_y = 2;
defparam syncreset_ctrl_X61_Y8.coord_z = 0;
defparam syncreset_ctrl_X61_Y8.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X61_Y9(
	.Din(),
	.Dout(SyncReset_X61_Y9_GND));
defparam syncreset_ctrl_X61_Y9.coord_x = 19;
defparam syncreset_ctrl_X61_Y9.coord_y = 7;
defparam syncreset_ctrl_X61_Y9.coord_z = 0;
defparam syncreset_ctrl_X61_Y9.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X62_Y1(
	.Din(),
	.Dout(SyncReset_X62_Y1_GND));
defparam syncreset_ctrl_X62_Y1.coord_x = 12;
defparam syncreset_ctrl_X62_Y1.coord_y = 1;
defparam syncreset_ctrl_X62_Y1.coord_z = 0;
defparam syncreset_ctrl_X62_Y1.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X62_Y10(
	.Din(),
	.Dout(SyncReset_X62_Y10_GND));
defparam syncreset_ctrl_X62_Y10.coord_x = 20;
defparam syncreset_ctrl_X62_Y10.coord_y = 12;
defparam syncreset_ctrl_X62_Y10.coord_z = 0;
defparam syncreset_ctrl_X62_Y10.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X62_Y11(
	.Din(),
	.Dout(SyncReset_X62_Y11_GND));
defparam syncreset_ctrl_X62_Y11.coord_x = 20;
defparam syncreset_ctrl_X62_Y11.coord_y = 9;
defparam syncreset_ctrl_X62_Y11.coord_z = 0;
defparam syncreset_ctrl_X62_Y11.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X62_Y2(
	.Din(),
	.Dout(SyncReset_X62_Y2_GND));
defparam syncreset_ctrl_X62_Y2.coord_x = 17;
defparam syncreset_ctrl_X62_Y2.coord_y = 6;
defparam syncreset_ctrl_X62_Y2.coord_z = 0;
defparam syncreset_ctrl_X62_Y2.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X62_Y3(
	.Din(),
	.Dout(SyncReset_X62_Y3_GND));
defparam syncreset_ctrl_X62_Y3.coord_x = 16;
defparam syncreset_ctrl_X62_Y3.coord_y = 6;
defparam syncreset_ctrl_X62_Y3.coord_z = 0;
defparam syncreset_ctrl_X62_Y3.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X62_Y4(
	.Din(),
	.Dout(SyncReset_X62_Y4_GND));
defparam syncreset_ctrl_X62_Y4.coord_x = 14;
defparam syncreset_ctrl_X62_Y4.coord_y = 3;
defparam syncreset_ctrl_X62_Y4.coord_z = 0;
defparam syncreset_ctrl_X62_Y4.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X62_Y5(
	.Din(),
	.Dout(SyncReset_X62_Y5_GND));
defparam syncreset_ctrl_X62_Y5.coord_x = 17;
defparam syncreset_ctrl_X62_Y5.coord_y = 10;
defparam syncreset_ctrl_X62_Y5.coord_z = 0;
defparam syncreset_ctrl_X62_Y5.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X62_Y6(
	.Din(),
	.Dout(SyncReset_X62_Y6_GND));
defparam syncreset_ctrl_X62_Y6.coord_x = 17;
defparam syncreset_ctrl_X62_Y6.coord_y = 12;
defparam syncreset_ctrl_X62_Y6.coord_z = 0;
defparam syncreset_ctrl_X62_Y6.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X62_Y7(
	.Din(),
	.Dout(SyncReset_X62_Y7_GND));
defparam syncreset_ctrl_X62_Y7.coord_x = 15;
defparam syncreset_ctrl_X62_Y7.coord_y = 6;
defparam syncreset_ctrl_X62_Y7.coord_z = 0;
defparam syncreset_ctrl_X62_Y7.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X62_Y8(
	.Din(),
	.Dout(SyncReset_X62_Y8_GND));
defparam syncreset_ctrl_X62_Y8.coord_x = 18;
defparam syncreset_ctrl_X62_Y8.coord_y = 2;
defparam syncreset_ctrl_X62_Y8.coord_z = 0;
defparam syncreset_ctrl_X62_Y8.SyncCtrlMux = 2'b00;

alta_syncctrl syncreset_ctrl_X62_Y9(
	.Din(),
	.Dout(SyncReset_X62_Y9_GND));
defparam syncreset_ctrl_X62_Y9.coord_x = 19;
defparam syncreset_ctrl_X62_Y9.coord_y = 11;
defparam syncreset_ctrl_X62_Y9.coord_z = 0;
defparam syncreset_ctrl_X62_Y9.SyncCtrlMux = 2'b00;

alta_slice sys_resetn(
	.A(vcc),
	.B(\rv32.resetn_out ),
	.C(vcc),
	.D(vcc),
	.Cin(),
	.Qin(),
	.Clk(),
	.AsyncReset(),
	.SyncReset(),
	.ShiftData(),
	.SyncLoad(),
	.LutOut(\sys_resetn~combout ),
	.Cout(),
	.Q());
defparam sys_resetn.coord_x = 20;
defparam sys_resetn.coord_y = 2;
defparam sys_resetn.coord_z = 4;
defparam sys_resetn.mask = 16'h3333;
defparam sys_resetn.modeMux = 1'b0;
defparam sys_resetn.FeedbackMux = 1'b0;
defparam sys_resetn.ShiftMux = 1'b0;
defparam sys_resetn.BypassEn = 1'b0;
defparam sys_resetn.CarryEnb = 1'b1;

alta_io_gclk \sys_resetn~clkctrl (
	.inclk(\sys_resetn~combout ),
	.outclk(\sys_resetn~clkctrl_outclk ));
defparam \sys_resetn~clkctrl .coord_x = 22;
defparam \sys_resetn~clkctrl .coord_y = 4;
defparam \sys_resetn~clkctrl .coord_z = 4;

endmodule
