module user_ip (
  input              CI_CK,
  input              CI_CS,
  input              CI_DAT,
  output tri0        CO_CK,
  output tri0        CO_CS,
  output tri0        CO_DAT,
  output tri0        D0,
  output tri0        D1,
  output tri0        D10,
  output tri0        D11,
  output tri0        D12,
  output tri0        D13,
  output tri0        D14,
  output tri0        D15,
  output tri0        D16,
  output tri0        D17,
  output tri0        D18,
  output tri0        D19,
  output tri0        D2,
  output tri0        D20,
  output tri0        D21,
  output tri0        D22,
  output tri0        D23,
  output tri0        D3,
  output tri0        D4,
  output tri0        D5,
  output tri0        D6,
  output tri0        D7,
  output tri0        D8,
  output tri0        D9,
  output tri0        LM_CK,
  input              LM_D0,
  input              LM_D1,
  input              LM_D2,
  input              LM_D3,
  input              LM_D4,
  input              LM_D5,
  output tri0        LM_LD,
  output tri0        SH1,
  output tri0        SH2,
  output tri0        SH3,
  output tri0        SH4,
  output tri0        SH5,
  output tri0        SH6,
  output tri0        ST1,
  output tri0        ST2,
  output tri0        csp_intr_in,
  input              sys_clock,
  input              bus_clock,
  input              resetn,
  input              stop,
  input       [1:0]  mem_ahb_htrans,
  input              mem_ahb_hready,
  input              mem_ahb_hwrite,
  input       [31:0] mem_ahb_haddr,
  input       [2:0]  mem_ahb_hsize,
  input       [2:0]  mem_ahb_hburst,
  input       [31:0] mem_ahb_hwdata,
  output tri1        mem_ahb_hreadyout,
  output tri0        mem_ahb_hresp,
  output tri0 [31:0] mem_ahb_hrdata,
  output tri0        slave_ahb_hsel,
  output tri1        slave_ahb_hready,
  input              slave_ahb_hreadyout,
  output tri0 [1:0]  slave_ahb_htrans,
  output tri0 [2:0]  slave_ahb_hsize,
  output tri0 [2:0]  slave_ahb_hburst,
  output tri0        slave_ahb_hwrite,
  output tri0 [31:0] slave_ahb_haddr,
  output tri0 [31:0] slave_ahb_hwdata,
  input              slave_ahb_hresp,
  input       [31:0] slave_ahb_hrdata,
  output tri0 [3:0]  ext_dma_DMACBREQ,
  output tri0 [3:0]  ext_dma_DMACLBREQ,
  output tri0 [3:0]  ext_dma_DMACSREQ,
  output tri0 [3:0]  ext_dma_DMACLSREQ,
  input       [3:0]  ext_dma_DMACCLR,
  input       [3:0]  ext_dma_DMACTC,
  output tri0 [3:0]  local_int
);
assign mem_ahb_hreadyout = 1'b1;
assign slave_ahb_hready  = 1'b1;
endmodule
